// nios_system.v

// Generated using ACDS version 12.1 177 at 2015.02.11.17:01:07

`timescale 1 ps / 1 ps
module nios_system (
		output wire [11:0] com_sdram_wire_addr,               //         com_sdram_wire.addr
		output wire [1:0]  com_sdram_wire_ba,                 //                       .ba
		output wire        com_sdram_wire_cas_n,              //                       .cas_n
		output wire        com_sdram_wire_cke,                //                       .cke
		output wire        com_sdram_wire_cs_n,               //                       .cs_n
		inout  wire [31:0] com_sdram_wire_dq,                 //                       .dq
		output wire [3:0]  com_sdram_wire_dqm,                //                       .dqm
		output wire        com_sdram_wire_ras_n,              //                       .ras_n
		output wire        com_sdram_wire_we_n,               //                       .we_n
		input  wire [3:0]  tse_conduit_connection_rgmii_in,   // tse_conduit_connection.rgmii_in
		output wire [3:0]  tse_conduit_connection_rgmii_out,  //                       .rgmii_out
		input  wire        tse_conduit_connection_rx_control, //                       .rx_control
		output wire        tse_conduit_connection_tx_control, //                       .tx_control
		input  wire        tse_conduit_connection_tx_clk,     //                       .tx_clk
		input  wire        tse_conduit_connection_rx_clk,     //                       .rx_clk
		input  wire        tse_conduit_connection_set_10,     //                       .set_10
		input  wire        tse_conduit_connection_set_1000,   //                       .set_1000
		output wire        tse_conduit_connection_ena_10,     //                       .ena_10
		output wire        tse_conduit_connection_eth_mode,   //                       .eth_mode
		output wire        tse_conduit_connection_mdio_out,   //                       .mdio_out
		output wire        tse_conduit_connection_mdio_oen,   //                       .mdio_oen
		input  wire        tse_conduit_connection_mdio_in,    //                       .mdio_in
		output wire        tse_conduit_connection_mdc,        //                       .mdc
		input  wire        reset_reset_n,                     //                  reset.reset_n
		input  wire        clk_clk                            //                    clk.clk
	);

	wire    [3:0] com_nios_instruction_master_burstcount;                                                                       // com_nios:i_burstcount -> com_nios_instruction_master_translator:av_burstcount
	wire          com_nios_instruction_master_waitrequest;                                                                      // com_nios_instruction_master_translator:av_waitrequest -> com_nios:i_waitrequest
	wire   [28:0] com_nios_instruction_master_address;                                                                          // com_nios:i_address -> com_nios_instruction_master_translator:av_address
	wire          com_nios_instruction_master_read;                                                                             // com_nios:i_read -> com_nios_instruction_master_translator:av_read
	wire   [31:0] com_nios_instruction_master_readdata;                                                                         // com_nios_instruction_master_translator:av_readdata -> com_nios:i_readdata
	wire          com_nios_instruction_master_readdatavalid;                                                                    // com_nios_instruction_master_translator:av_readdatavalid -> com_nios:i_readdatavalid
	wire    [3:0] com_nios_data_master_burstcount;                                                                              // com_nios:d_burstcount -> com_nios_data_master_translator:av_burstcount
	wire          com_nios_data_master_waitrequest;                                                                             // com_nios_data_master_translator:av_waitrequest -> com_nios:d_waitrequest
	wire   [31:0] com_nios_data_master_writedata;                                                                               // com_nios:d_writedata -> com_nios_data_master_translator:av_writedata
	wire   [28:0] com_nios_data_master_address;                                                                                 // com_nios:d_address -> com_nios_data_master_translator:av_address
	wire          com_nios_data_master_write;                                                                                   // com_nios:d_write -> com_nios_data_master_translator:av_write
	wire          com_nios_data_master_read;                                                                                    // com_nios:d_read -> com_nios_data_master_translator:av_read
	wire   [31:0] com_nios_data_master_readdata;                                                                                // com_nios_data_master_translator:av_readdata -> com_nios:d_readdata
	wire          com_nios_data_master_debugaccess;                                                                             // com_nios:jtag_debug_module_debugaccess_to_roms -> com_nios_data_master_translator:av_debugaccess
	wire          com_nios_data_master_readdatavalid;                                                                           // com_nios_data_master_translator:av_readdatavalid -> com_nios:d_readdatavalid
	wire    [3:0] com_nios_data_master_byteenable;                                                                              // com_nios:d_byteenable -> com_nios_data_master_translator:av_byteenable
	wire          carcontrol_nios_data_master_waitrequest;                                                                      // carControl_nios_data_master_translator:av_waitrequest -> carControl_nios:d_waitrequest
	wire   [31:0] carcontrol_nios_data_master_writedata;                                                                        // carControl_nios:d_writedata -> carControl_nios_data_master_translator:av_writedata
	wire   [28:0] carcontrol_nios_data_master_address;                                                                          // carControl_nios:d_address -> carControl_nios_data_master_translator:av_address
	wire          carcontrol_nios_data_master_write;                                                                            // carControl_nios:d_write -> carControl_nios_data_master_translator:av_write
	wire          carcontrol_nios_data_master_read;                                                                             // carControl_nios:d_read -> carControl_nios_data_master_translator:av_read
	wire   [31:0] carcontrol_nios_data_master_readdata;                                                                         // carControl_nios_data_master_translator:av_readdata -> carControl_nios:d_readdata
	wire          carcontrol_nios_data_master_debugaccess;                                                                      // carControl_nios:jtag_debug_module_debugaccess_to_roms -> carControl_nios_data_master_translator:av_debugaccess
	wire    [3:0] carcontrol_nios_data_master_byteenable;                                                                       // carControl_nios:d_byteenable -> carControl_nios_data_master_translator:av_byteenable
	wire          carcontrol_nios_instruction_master_waitrequest;                                                               // carControl_nios_instruction_master_translator:av_waitrequest -> carControl_nios:i_waitrequest
	wire   [28:0] carcontrol_nios_instruction_master_address;                                                                   // carControl_nios:i_address -> carControl_nios_instruction_master_translator:av_address
	wire          carcontrol_nios_instruction_master_read;                                                                      // carControl_nios:i_read -> carControl_nios_instruction_master_translator:av_read
	wire   [31:0] carcontrol_nios_instruction_master_readdata;                                                                  // carControl_nios_instruction_master_translator:av_readdata -> carControl_nios:i_readdata
	wire          carcontrol_nios_instruction_master_readdatavalid;                                                             // carControl_nios_instruction_master_translator:av_readdatavalid -> carControl_nios:i_readdatavalid
	wire          ethernet_subsystem_sgdma_rx_m_write_waitrequest;                                                              // ethernet_subsystem_sgdma_rx_m_write_translator:av_waitrequest -> ethernet_subsystem:sgdma_rx_m_write_waitrequest
	wire   [31:0] ethernet_subsystem_sgdma_rx_m_write_writedata;                                                                // ethernet_subsystem:sgdma_rx_m_write_writedata -> ethernet_subsystem_sgdma_rx_m_write_translator:av_writedata
	wire   [31:0] ethernet_subsystem_sgdma_rx_m_write_address;                                                                  // ethernet_subsystem:sgdma_rx_m_write_address -> ethernet_subsystem_sgdma_rx_m_write_translator:av_address
	wire          ethernet_subsystem_sgdma_rx_m_write_write;                                                                    // ethernet_subsystem:sgdma_rx_m_write_write -> ethernet_subsystem_sgdma_rx_m_write_translator:av_write
	wire    [3:0] ethernet_subsystem_sgdma_rx_m_write_byteenable;                                                               // ethernet_subsystem:sgdma_rx_m_write_byteenable -> ethernet_subsystem_sgdma_rx_m_write_translator:av_byteenable
	wire          ethernet_subsystem_sgdma_tx_m_read_waitrequest;                                                               // ethernet_subsystem_sgdma_tx_m_read_translator:av_waitrequest -> ethernet_subsystem:sgdma_tx_m_read_waitrequest
	wire   [31:0] ethernet_subsystem_sgdma_tx_m_read_address;                                                                   // ethernet_subsystem:sgdma_tx_m_read_address -> ethernet_subsystem_sgdma_tx_m_read_translator:av_address
	wire          ethernet_subsystem_sgdma_tx_m_read_read;                                                                      // ethernet_subsystem:sgdma_tx_m_read_read -> ethernet_subsystem_sgdma_tx_m_read_translator:av_read
	wire   [31:0] ethernet_subsystem_sgdma_tx_m_read_readdata;                                                                  // ethernet_subsystem_sgdma_tx_m_read_translator:av_readdata -> ethernet_subsystem:sgdma_tx_m_read_readdata
	wire          ethernet_subsystem_sgdma_tx_m_read_readdatavalid;                                                             // ethernet_subsystem_sgdma_tx_m_read_translator:av_readdatavalid -> ethernet_subsystem:sgdma_tx_m_read_readdatavalid
	wire   [31:0] com_nios_jtag_debug_module_translator_avalon_anti_slave_0_writedata;                                          // com_nios_jtag_debug_module_translator:av_writedata -> com_nios:jtag_debug_module_writedata
	wire    [8:0] com_nios_jtag_debug_module_translator_avalon_anti_slave_0_address;                                            // com_nios_jtag_debug_module_translator:av_address -> com_nios:jtag_debug_module_address
	wire          com_nios_jtag_debug_module_translator_avalon_anti_slave_0_chipselect;                                         // com_nios_jtag_debug_module_translator:av_chipselect -> com_nios:jtag_debug_module_select
	wire          com_nios_jtag_debug_module_translator_avalon_anti_slave_0_write;                                              // com_nios_jtag_debug_module_translator:av_write -> com_nios:jtag_debug_module_write
	wire   [31:0] com_nios_jtag_debug_module_translator_avalon_anti_slave_0_readdata;                                           // com_nios:jtag_debug_module_readdata -> com_nios_jtag_debug_module_translator:av_readdata
	wire          com_nios_jtag_debug_module_translator_avalon_anti_slave_0_begintransfer;                                      // com_nios_jtag_debug_module_translator:av_begintransfer -> com_nios:jtag_debug_module_begintransfer
	wire          com_nios_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess;                                        // com_nios_jtag_debug_module_translator:av_debugaccess -> com_nios:jtag_debug_module_debugaccess
	wire    [3:0] com_nios_jtag_debug_module_translator_avalon_anti_slave_0_byteenable;                                         // com_nios_jtag_debug_module_translator:av_byteenable -> com_nios:jtag_debug_module_byteenable
	wire          com_memory_s1_translator_avalon_anti_slave_0_waitrequest;                                                     // com_memory:za_waitrequest -> com_memory_s1_translator:av_waitrequest
	wire   [31:0] com_memory_s1_translator_avalon_anti_slave_0_writedata;                                                       // com_memory_s1_translator:av_writedata -> com_memory:az_data
	wire   [23:0] com_memory_s1_translator_avalon_anti_slave_0_address;                                                         // com_memory_s1_translator:av_address -> com_memory:az_addr
	wire          com_memory_s1_translator_avalon_anti_slave_0_chipselect;                                                      // com_memory_s1_translator:av_chipselect -> com_memory:az_cs
	wire          com_memory_s1_translator_avalon_anti_slave_0_write;                                                           // com_memory_s1_translator:av_write -> com_memory:az_wr_n
	wire          com_memory_s1_translator_avalon_anti_slave_0_read;                                                            // com_memory_s1_translator:av_read -> com_memory:az_rd_n
	wire   [31:0] com_memory_s1_translator_avalon_anti_slave_0_readdata;                                                        // com_memory:za_data -> com_memory_s1_translator:av_readdata
	wire          com_memory_s1_translator_avalon_anti_slave_0_readdatavalid;                                                   // com_memory:za_valid -> com_memory_s1_translator:av_readdatavalid
	wire    [3:0] com_memory_s1_translator_avalon_anti_slave_0_byteenable;                                                      // com_memory_s1_translator:av_byteenable -> com_memory:az_be_n
	wire          jtaguart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest;                                      // jtaguart_0:av_waitrequest -> jtaguart_0_avalon_jtag_slave_translator:av_waitrequest
	wire   [31:0] jtaguart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata;                                        // jtaguart_0_avalon_jtag_slave_translator:av_writedata -> jtaguart_0:av_writedata
	wire    [0:0] jtaguart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_address;                                          // jtaguart_0_avalon_jtag_slave_translator:av_address -> jtaguart_0:av_address
	wire          jtaguart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect;                                       // jtaguart_0_avalon_jtag_slave_translator:av_chipselect -> jtaguart_0:av_chipselect
	wire          jtaguart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_write;                                            // jtaguart_0_avalon_jtag_slave_translator:av_write -> jtaguart_0:av_write_n
	wire          jtaguart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_read;                                             // jtaguart_0_avalon_jtag_slave_translator:av_read -> jtaguart_0:av_read_n
	wire   [31:0] jtaguart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata;                                         // jtaguart_0:av_readdata -> jtaguart_0_avalon_jtag_slave_translator:av_readdata
	wire   [31:0] shared_memory_mutex_s1_translator_avalon_anti_slave_0_writedata;                                              // shared_memory_mutex_s1_translator:av_writedata -> shared_memory_mutex:data_from_cpu
	wire    [0:0] shared_memory_mutex_s1_translator_avalon_anti_slave_0_address;                                                // shared_memory_mutex_s1_translator:av_address -> shared_memory_mutex:address
	wire          shared_memory_mutex_s1_translator_avalon_anti_slave_0_chipselect;                                             // shared_memory_mutex_s1_translator:av_chipselect -> shared_memory_mutex:chipselect
	wire          shared_memory_mutex_s1_translator_avalon_anti_slave_0_write;                                                  // shared_memory_mutex_s1_translator:av_write -> shared_memory_mutex:write
	wire          shared_memory_mutex_s1_translator_avalon_anti_slave_0_read;                                                   // shared_memory_mutex_s1_translator:av_read -> shared_memory_mutex:read
	wire   [31:0] shared_memory_mutex_s1_translator_avalon_anti_slave_0_readdata;                                               // shared_memory_mutex:data_to_cpu -> shared_memory_mutex_s1_translator:av_readdata
	wire   [15:0] com_timer_s1_translator_avalon_anti_slave_0_writedata;                                                        // com_timer_s1_translator:av_writedata -> com_timer:writedata
	wire    [2:0] com_timer_s1_translator_avalon_anti_slave_0_address;                                                          // com_timer_s1_translator:av_address -> com_timer:address
	wire          com_timer_s1_translator_avalon_anti_slave_0_chipselect;                                                       // com_timer_s1_translator:av_chipselect -> com_timer:chipselect
	wire          com_timer_s1_translator_avalon_anti_slave_0_write;                                                            // com_timer_s1_translator:av_write -> com_timer:write_n
	wire   [15:0] com_timer_s1_translator_avalon_anti_slave_0_readdata;                                                         // com_timer:readdata -> com_timer_s1_translator:av_readdata
	wire          ethernet_subsystem_ethernet_bridge_s0_translator_avalon_anti_slave_0_waitrequest;                             // ethernet_subsystem:ethernet_bridge_s0_waitrequest -> ethernet_subsystem_ethernet_bridge_s0_translator:av_waitrequest
	wire    [0:0] ethernet_subsystem_ethernet_bridge_s0_translator_avalon_anti_slave_0_burstcount;                              // ethernet_subsystem_ethernet_bridge_s0_translator:av_burstcount -> ethernet_subsystem:ethernet_bridge_s0_burstcount
	wire   [31:0] ethernet_subsystem_ethernet_bridge_s0_translator_avalon_anti_slave_0_writedata;                               // ethernet_subsystem_ethernet_bridge_s0_translator:av_writedata -> ethernet_subsystem:ethernet_bridge_s0_writedata
	wire   [10:0] ethernet_subsystem_ethernet_bridge_s0_translator_avalon_anti_slave_0_address;                                 // ethernet_subsystem_ethernet_bridge_s0_translator:av_address -> ethernet_subsystem:ethernet_bridge_s0_address
	wire          ethernet_subsystem_ethernet_bridge_s0_translator_avalon_anti_slave_0_write;                                   // ethernet_subsystem_ethernet_bridge_s0_translator:av_write -> ethernet_subsystem:ethernet_bridge_s0_write
	wire          ethernet_subsystem_ethernet_bridge_s0_translator_avalon_anti_slave_0_read;                                    // ethernet_subsystem_ethernet_bridge_s0_translator:av_read -> ethernet_subsystem:ethernet_bridge_s0_read
	wire   [31:0] ethernet_subsystem_ethernet_bridge_s0_translator_avalon_anti_slave_0_readdata;                                // ethernet_subsystem:ethernet_bridge_s0_readdata -> ethernet_subsystem_ethernet_bridge_s0_translator:av_readdata
	wire          ethernet_subsystem_ethernet_bridge_s0_translator_avalon_anti_slave_0_debugaccess;                             // ethernet_subsystem_ethernet_bridge_s0_translator:av_debugaccess -> ethernet_subsystem:ethernet_bridge_s0_debugaccess
	wire          ethernet_subsystem_ethernet_bridge_s0_translator_avalon_anti_slave_0_readdatavalid;                           // ethernet_subsystem:ethernet_bridge_s0_readdatavalid -> ethernet_subsystem_ethernet_bridge_s0_translator:av_readdatavalid
	wire    [3:0] ethernet_subsystem_ethernet_bridge_s0_translator_avalon_anti_slave_0_byteenable;                              // ethernet_subsystem_ethernet_bridge_s0_translator:av_byteenable -> ethernet_subsystem:ethernet_bridge_s0_byteenable
	wire   [31:0] ethernet_subsystem_descriptor_memory_s2_translator_avalon_anti_slave_0_writedata;                             // ethernet_subsystem_descriptor_memory_s2_translator:av_writedata -> ethernet_subsystem:descriptor_memory_s2_writedata
	wire   [10:0] ethernet_subsystem_descriptor_memory_s2_translator_avalon_anti_slave_0_address;                               // ethernet_subsystem_descriptor_memory_s2_translator:av_address -> ethernet_subsystem:descriptor_memory_s2_address
	wire          ethernet_subsystem_descriptor_memory_s2_translator_avalon_anti_slave_0_chipselect;                            // ethernet_subsystem_descriptor_memory_s2_translator:av_chipselect -> ethernet_subsystem:descriptor_memory_s2_chipselect
	wire          ethernet_subsystem_descriptor_memory_s2_translator_avalon_anti_slave_0_clken;                                 // ethernet_subsystem_descriptor_memory_s2_translator:av_clken -> ethernet_subsystem:descriptor_memory_s2_clken
	wire          ethernet_subsystem_descriptor_memory_s2_translator_avalon_anti_slave_0_write;                                 // ethernet_subsystem_descriptor_memory_s2_translator:av_write -> ethernet_subsystem:descriptor_memory_s2_write
	wire   [31:0] ethernet_subsystem_descriptor_memory_s2_translator_avalon_anti_slave_0_readdata;                              // ethernet_subsystem:descriptor_memory_s2_readdata -> ethernet_subsystem_descriptor_memory_s2_translator:av_readdata
	wire    [3:0] ethernet_subsystem_descriptor_memory_s2_translator_avalon_anti_slave_0_byteenable;                            // ethernet_subsystem_descriptor_memory_s2_translator:av_byteenable -> ethernet_subsystem:descriptor_memory_s2_byteenable
	wire          prio_arbiter_0_s0_translator_avalon_anti_slave_0_waitrequest;                                                 // prio_arbiter_0:AVS_S0_WAITREQUEST -> prio_arbiter_0_s0_translator:av_waitrequest
	wire   [31:0] prio_arbiter_0_s0_translator_avalon_anti_slave_0_writedata;                                                   // prio_arbiter_0_s0_translator:av_writedata -> prio_arbiter_0:AVS_S0_WRITEDATA
	wire   [25:0] prio_arbiter_0_s0_translator_avalon_anti_slave_0_address;                                                     // prio_arbiter_0_s0_translator:av_address -> prio_arbiter_0:AVS_S0_ADDRESS
	wire          prio_arbiter_0_s0_translator_avalon_anti_slave_0_chipselect;                                                  // prio_arbiter_0_s0_translator:av_chipselect -> prio_arbiter_0:AVS_S0_CHIPSELECT
	wire          prio_arbiter_0_s0_translator_avalon_anti_slave_0_write;                                                       // prio_arbiter_0_s0_translator:av_write -> prio_arbiter_0:AVS_S0_WRITE
	wire          prio_arbiter_0_s0_translator_avalon_anti_slave_0_read;                                                        // prio_arbiter_0_s0_translator:av_read -> prio_arbiter_0:AVS_S0_READ
	wire   [31:0] prio_arbiter_0_s0_translator_avalon_anti_slave_0_readdata;                                                    // prio_arbiter_0:AVS_S0_READDATA -> prio_arbiter_0_s0_translator:av_readdata
	wire          prio_arbiter_0_s0_translator_avalon_anti_slave_0_readdatavalid;                                               // prio_arbiter_0:AVS_S0_READDATAVALID -> prio_arbiter_0_s0_translator:av_readdatavalid
	wire    [3:0] prio_arbiter_0_s0_translator_avalon_anti_slave_0_byteenable;                                                  // prio_arbiter_0_s0_translator:av_byteenable -> prio_arbiter_0:AVS_S0_BYTEENABLE
	wire   [31:0] carcontrol_nios_jtag_debug_module_translator_avalon_anti_slave_0_writedata;                                   // carControl_nios_jtag_debug_module_translator:av_writedata -> carControl_nios:jtag_debug_module_writedata
	wire    [8:0] carcontrol_nios_jtag_debug_module_translator_avalon_anti_slave_0_address;                                     // carControl_nios_jtag_debug_module_translator:av_address -> carControl_nios:jtag_debug_module_address
	wire          carcontrol_nios_jtag_debug_module_translator_avalon_anti_slave_0_chipselect;                                  // carControl_nios_jtag_debug_module_translator:av_chipselect -> carControl_nios:jtag_debug_module_select
	wire          carcontrol_nios_jtag_debug_module_translator_avalon_anti_slave_0_write;                                       // carControl_nios_jtag_debug_module_translator:av_write -> carControl_nios:jtag_debug_module_write
	wire   [31:0] carcontrol_nios_jtag_debug_module_translator_avalon_anti_slave_0_readdata;                                    // carControl_nios:jtag_debug_module_readdata -> carControl_nios_jtag_debug_module_translator:av_readdata
	wire          carcontrol_nios_jtag_debug_module_translator_avalon_anti_slave_0_begintransfer;                               // carControl_nios_jtag_debug_module_translator:av_begintransfer -> carControl_nios:jtag_debug_module_begintransfer
	wire          carcontrol_nios_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess;                                 // carControl_nios_jtag_debug_module_translator:av_debugaccess -> carControl_nios:jtag_debug_module_debugaccess
	wire    [3:0] carcontrol_nios_jtag_debug_module_translator_avalon_anti_slave_0_byteenable;                                  // carControl_nios_jtag_debug_module_translator:av_byteenable -> carControl_nios:jtag_debug_module_byteenable
	wire   [31:0] onchip_memory2_0_s1_translator_avalon_anti_slave_0_writedata;                                                 // onchip_memory2_0_s1_translator:av_writedata -> onchip_memory2_0:writedata
	wire   [15:0] onchip_memory2_0_s1_translator_avalon_anti_slave_0_address;                                                   // onchip_memory2_0_s1_translator:av_address -> onchip_memory2_0:address
	wire          onchip_memory2_0_s1_translator_avalon_anti_slave_0_chipselect;                                                // onchip_memory2_0_s1_translator:av_chipselect -> onchip_memory2_0:chipselect
	wire          onchip_memory2_0_s1_translator_avalon_anti_slave_0_clken;                                                     // onchip_memory2_0_s1_translator:av_clken -> onchip_memory2_0:clken
	wire          onchip_memory2_0_s1_translator_avalon_anti_slave_0_write;                                                     // onchip_memory2_0_s1_translator:av_write -> onchip_memory2_0:write
	wire   [31:0] onchip_memory2_0_s1_translator_avalon_anti_slave_0_readdata;                                                  // onchip_memory2_0:readdata -> onchip_memory2_0_s1_translator:av_readdata
	wire    [3:0] onchip_memory2_0_s1_translator_avalon_anti_slave_0_byteenable;                                                // onchip_memory2_0_s1_translator:av_byteenable -> onchip_memory2_0:byteenable
	wire          jtaguart_1_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest;                                      // jtaguart_1:av_waitrequest -> jtaguart_1_avalon_jtag_slave_translator:av_waitrequest
	wire   [31:0] jtaguart_1_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata;                                        // jtaguart_1_avalon_jtag_slave_translator:av_writedata -> jtaguart_1:av_writedata
	wire    [0:0] jtaguart_1_avalon_jtag_slave_translator_avalon_anti_slave_0_address;                                          // jtaguart_1_avalon_jtag_slave_translator:av_address -> jtaguart_1:av_address
	wire          jtaguart_1_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect;                                       // jtaguart_1_avalon_jtag_slave_translator:av_chipselect -> jtaguart_1:av_chipselect
	wire          jtaguart_1_avalon_jtag_slave_translator_avalon_anti_slave_0_write;                                            // jtaguart_1_avalon_jtag_slave_translator:av_write -> jtaguart_1:av_write_n
	wire          jtaguart_1_avalon_jtag_slave_translator_avalon_anti_slave_0_read;                                             // jtaguart_1_avalon_jtag_slave_translator:av_read -> jtaguart_1:av_read_n
	wire   [31:0] jtaguart_1_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata;                                         // jtaguart_1:av_readdata -> jtaguart_1_avalon_jtag_slave_translator:av_readdata
	wire          prio_arbiter_0_s1_translator_avalon_anti_slave_0_waitrequest;                                                 // prio_arbiter_0:AVS_S1_WAITREQUEST -> prio_arbiter_0_s1_translator:av_waitrequest
	wire   [31:0] prio_arbiter_0_s1_translator_avalon_anti_slave_0_writedata;                                                   // prio_arbiter_0_s1_translator:av_writedata -> prio_arbiter_0:AVS_S1_WRITEDATA
	wire   [25:0] prio_arbiter_0_s1_translator_avalon_anti_slave_0_address;                                                     // prio_arbiter_0_s1_translator:av_address -> prio_arbiter_0:AVS_S1_ADDRESS
	wire          prio_arbiter_0_s1_translator_avalon_anti_slave_0_chipselect;                                                  // prio_arbiter_0_s1_translator:av_chipselect -> prio_arbiter_0:AVS_S1_CHIPSELECT
	wire          prio_arbiter_0_s1_translator_avalon_anti_slave_0_write;                                                       // prio_arbiter_0_s1_translator:av_write -> prio_arbiter_0:AVS_S1_WRITE
	wire          prio_arbiter_0_s1_translator_avalon_anti_slave_0_read;                                                        // prio_arbiter_0_s1_translator:av_read -> prio_arbiter_0:AVS_S1_READ
	wire   [31:0] prio_arbiter_0_s1_translator_avalon_anti_slave_0_readdata;                                                    // prio_arbiter_0:AVS_S1_READDATA -> prio_arbiter_0_s1_translator:av_readdata
	wire          prio_arbiter_0_s1_translator_avalon_anti_slave_0_readdatavalid;                                               // prio_arbiter_0:AVS_S1_READDATAVALID -> prio_arbiter_0_s1_translator:av_readdatavalid
	wire    [3:0] prio_arbiter_0_s1_translator_avalon_anti_slave_0_byteenable;                                                  // prio_arbiter_0_s1_translator:av_byteenable -> prio_arbiter_0:AVS_S1_BYTEENABLE
	wire          prio_arbiter_0_m1_waitrequest;                                                                                // prio_arbiter_0_m1_translator:av_waitrequest -> prio_arbiter_0:AVM_M1_WAITREQUEST
	wire   [31:0] prio_arbiter_0_m1_writedata;                                                                                  // prio_arbiter_0:AVM_M1_WRITEDATA -> prio_arbiter_0_m1_translator:av_writedata
	wire   [27:0] prio_arbiter_0_m1_address;                                                                                    // prio_arbiter_0:AVM_M1_ADDRESS -> prio_arbiter_0_m1_translator:av_address
	wire          prio_arbiter_0_m1_write;                                                                                      // prio_arbiter_0:AVM_M1_WRITE -> prio_arbiter_0_m1_translator:av_write
	wire          prio_arbiter_0_m1_read;                                                                                       // prio_arbiter_0:AVM_M1_READ -> prio_arbiter_0_m1_translator:av_read
	wire   [31:0] prio_arbiter_0_m1_readdata;                                                                                   // prio_arbiter_0_m1_translator:av_readdata -> prio_arbiter_0:AVM_M1_READDATA
	wire          prio_arbiter_0_m1_readdatavalid;                                                                              // prio_arbiter_0_m1_translator:av_readdatavalid -> prio_arbiter_0:AVM_M1_READDATAVALID
	wire    [3:0] prio_arbiter_0_m1_byteenable;                                                                                 // prio_arbiter_0:AVM_M1_BYTEENABLE -> prio_arbiter_0_m1_translator:av_byteenable
	wire          prio_arbiter_0_m1_translator_avalon_universal_master_0_waitrequest;                                           // shared_memory_s1_translator:uav_waitrequest -> prio_arbiter_0_m1_translator:uav_waitrequest
	wire    [2:0] prio_arbiter_0_m1_translator_avalon_universal_master_0_burstcount;                                            // prio_arbiter_0_m1_translator:uav_burstcount -> shared_memory_s1_translator:uav_burstcount
	wire   [31:0] prio_arbiter_0_m1_translator_avalon_universal_master_0_writedata;                                             // prio_arbiter_0_m1_translator:uav_writedata -> shared_memory_s1_translator:uav_writedata
	wire   [27:0] prio_arbiter_0_m1_translator_avalon_universal_master_0_address;                                               // prio_arbiter_0_m1_translator:uav_address -> shared_memory_s1_translator:uav_address
	wire          prio_arbiter_0_m1_translator_avalon_universal_master_0_lock;                                                  // prio_arbiter_0_m1_translator:uav_lock -> shared_memory_s1_translator:uav_lock
	wire          prio_arbiter_0_m1_translator_avalon_universal_master_0_write;                                                 // prio_arbiter_0_m1_translator:uav_write -> shared_memory_s1_translator:uav_write
	wire          prio_arbiter_0_m1_translator_avalon_universal_master_0_read;                                                  // prio_arbiter_0_m1_translator:uav_read -> shared_memory_s1_translator:uav_read
	wire   [31:0] prio_arbiter_0_m1_translator_avalon_universal_master_0_readdata;                                              // shared_memory_s1_translator:uav_readdata -> prio_arbiter_0_m1_translator:uav_readdata
	wire          prio_arbiter_0_m1_translator_avalon_universal_master_0_debugaccess;                                           // prio_arbiter_0_m1_translator:uav_debugaccess -> shared_memory_s1_translator:uav_debugaccess
	wire    [3:0] prio_arbiter_0_m1_translator_avalon_universal_master_0_byteenable;                                            // prio_arbiter_0_m1_translator:uav_byteenable -> shared_memory_s1_translator:uav_byteenable
	wire          prio_arbiter_0_m1_translator_avalon_universal_master_0_readdatavalid;                                         // shared_memory_s1_translator:uav_readdatavalid -> prio_arbiter_0_m1_translator:uav_readdatavalid
	wire   [31:0] shared_memory_s1_translator_avalon_anti_slave_0_writedata;                                                    // shared_memory_s1_translator:av_writedata -> shared_memory:writedata
	wire    [9:0] shared_memory_s1_translator_avalon_anti_slave_0_address;                                                      // shared_memory_s1_translator:av_address -> shared_memory:address
	wire          shared_memory_s1_translator_avalon_anti_slave_0_chipselect;                                                   // shared_memory_s1_translator:av_chipselect -> shared_memory:chipselect
	wire          shared_memory_s1_translator_avalon_anti_slave_0_clken;                                                        // shared_memory_s1_translator:av_clken -> shared_memory:clken
	wire          shared_memory_s1_translator_avalon_anti_slave_0_write;                                                        // shared_memory_s1_translator:av_write -> shared_memory:write
	wire   [31:0] shared_memory_s1_translator_avalon_anti_slave_0_readdata;                                                     // shared_memory:readdata -> shared_memory_s1_translator:av_readdata
	wire    [3:0] shared_memory_s1_translator_avalon_anti_slave_0_byteenable;                                                   // shared_memory_s1_translator:av_byteenable -> shared_memory:byteenable
	wire    [3:0] traffic_gen_0_avalon_master_0_burstcount;                                                                     // traffic_gen_0:MASTER_BURSTCOUNT_AVM -> traffic_gen_0_avalon_master_0_translator:av_burstcount
	wire          traffic_gen_0_avalon_master_0_waitrequest;                                                                    // traffic_gen_0_avalon_master_0_translator:av_waitrequest -> traffic_gen_0:MASTER_WAITREQUEST_AVM
	wire   [31:0] traffic_gen_0_avalon_master_0_writedata;                                                                      // traffic_gen_0:MASTER_WRITEDATA_AVM -> traffic_gen_0_avalon_master_0_translator:av_writedata
	wire   [27:0] traffic_gen_0_avalon_master_0_address;                                                                        // traffic_gen_0:MASTER_ADDRES_AVM -> traffic_gen_0_avalon_master_0_translator:av_address
	wire          traffic_gen_0_avalon_master_0_write;                                                                          // traffic_gen_0:MASTER_WRITE_AVM -> traffic_gen_0_avalon_master_0_translator:av_write
	wire          traffic_gen_0_avalon_master_0_read;                                                                           // traffic_gen_0:MASTER_READ_AVM -> traffic_gen_0_avalon_master_0_translator:av_read
	wire   [31:0] traffic_gen_0_avalon_master_0_readdata;                                                                       // traffic_gen_0_avalon_master_0_translator:av_readdata -> traffic_gen_0:MASTER_READ_DATA_AVM
	wire          traffic_gen_0_avalon_master_0_readdatavalid;                                                                  // traffic_gen_0_avalon_master_0_translator:av_readdatavalid -> traffic_gen_0:MASTER_READDATAVALID_AVM
	wire    [3:0] traffic_gen_0_avalon_master_0_byteenable;                                                                     // traffic_gen_0:MASTER_BYTEENABLE_AVM -> traffic_gen_0_avalon_master_0_translator:av_byteenable
	wire          prio_arbiter_0_s2_translator_avalon_anti_slave_0_waitrequest;                                                 // prio_arbiter_0:AVS_S2_WAITREQUEST -> prio_arbiter_0_s2_translator:av_waitrequest
	wire   [31:0] prio_arbiter_0_s2_translator_avalon_anti_slave_0_writedata;                                                   // prio_arbiter_0_s2_translator:av_writedata -> prio_arbiter_0:AVS_S2_WRITEDATA
	wire   [25:0] prio_arbiter_0_s2_translator_avalon_anti_slave_0_address;                                                     // prio_arbiter_0_s2_translator:av_address -> prio_arbiter_0:AVS_S2_ADDRESS
	wire          prio_arbiter_0_s2_translator_avalon_anti_slave_0_chipselect;                                                  // prio_arbiter_0_s2_translator:av_chipselect -> prio_arbiter_0:AVS_S2_CHIPSELECT
	wire          prio_arbiter_0_s2_translator_avalon_anti_slave_0_write;                                                       // prio_arbiter_0_s2_translator:av_write -> prio_arbiter_0:AVS_S2_WRITE
	wire          prio_arbiter_0_s2_translator_avalon_anti_slave_0_read;                                                        // prio_arbiter_0_s2_translator:av_read -> prio_arbiter_0:AVS_S2_READ
	wire   [31:0] prio_arbiter_0_s2_translator_avalon_anti_slave_0_readdata;                                                    // prio_arbiter_0:AVS_S2_READDATA -> prio_arbiter_0_s2_translator:av_readdata
	wire          prio_arbiter_0_s2_translator_avalon_anti_slave_0_readdatavalid;                                               // prio_arbiter_0:AVS_S2_READDATAVALID -> prio_arbiter_0_s2_translator:av_readdatavalid
	wire    [3:0] prio_arbiter_0_s2_translator_avalon_anti_slave_0_byteenable;                                                  // prio_arbiter_0_s2_translator:av_byteenable -> prio_arbiter_0:AVS_S2_BYTEENABLE
	wire    [3:0] traffic_gen_1_avalon_master_0_burstcount;                                                                     // traffic_gen_1:MASTER_BURSTCOUNT_AVM -> traffic_gen_1_avalon_master_0_translator:av_burstcount
	wire          traffic_gen_1_avalon_master_0_waitrequest;                                                                    // traffic_gen_1_avalon_master_0_translator:av_waitrequest -> traffic_gen_1:MASTER_WAITREQUEST_AVM
	wire   [31:0] traffic_gen_1_avalon_master_0_writedata;                                                                      // traffic_gen_1:MASTER_WRITEDATA_AVM -> traffic_gen_1_avalon_master_0_translator:av_writedata
	wire   [27:0] traffic_gen_1_avalon_master_0_address;                                                                        // traffic_gen_1:MASTER_ADDRES_AVM -> traffic_gen_1_avalon_master_0_translator:av_address
	wire          traffic_gen_1_avalon_master_0_write;                                                                          // traffic_gen_1:MASTER_WRITE_AVM -> traffic_gen_1_avalon_master_0_translator:av_write
	wire          traffic_gen_1_avalon_master_0_read;                                                                           // traffic_gen_1:MASTER_READ_AVM -> traffic_gen_1_avalon_master_0_translator:av_read
	wire   [31:0] traffic_gen_1_avalon_master_0_readdata;                                                                       // traffic_gen_1_avalon_master_0_translator:av_readdata -> traffic_gen_1:MASTER_READ_DATA_AVM
	wire          traffic_gen_1_avalon_master_0_readdatavalid;                                                                  // traffic_gen_1_avalon_master_0_translator:av_readdatavalid -> traffic_gen_1:MASTER_READDATAVALID_AVM
	wire    [3:0] traffic_gen_1_avalon_master_0_byteenable;                                                                     // traffic_gen_1:MASTER_BYTEENABLE_AVM -> traffic_gen_1_avalon_master_0_translator:av_byteenable
	wire          prio_arbiter_0_s3_translator_avalon_anti_slave_0_waitrequest;                                                 // prio_arbiter_0:AVS_S3_WAITREQUEST -> prio_arbiter_0_s3_translator:av_waitrequest
	wire   [31:0] prio_arbiter_0_s3_translator_avalon_anti_slave_0_writedata;                                                   // prio_arbiter_0_s3_translator:av_writedata -> prio_arbiter_0:AVS_S3_WRITEDATA
	wire   [25:0] prio_arbiter_0_s3_translator_avalon_anti_slave_0_address;                                                     // prio_arbiter_0_s3_translator:av_address -> prio_arbiter_0:AVS_S3_ADDRESS
	wire          prio_arbiter_0_s3_translator_avalon_anti_slave_0_chipselect;                                                  // prio_arbiter_0_s3_translator:av_chipselect -> prio_arbiter_0:AVS_S3_CHIPSELECT
	wire          prio_arbiter_0_s3_translator_avalon_anti_slave_0_write;                                                       // prio_arbiter_0_s3_translator:av_write -> prio_arbiter_0:AVS_S3_WRITE
	wire          prio_arbiter_0_s3_translator_avalon_anti_slave_0_read;                                                        // prio_arbiter_0_s3_translator:av_read -> prio_arbiter_0:AVS_S3_READ
	wire   [31:0] prio_arbiter_0_s3_translator_avalon_anti_slave_0_readdata;                                                    // prio_arbiter_0:AVS_S3_READDATA -> prio_arbiter_0_s3_translator:av_readdata
	wire          prio_arbiter_0_s3_translator_avalon_anti_slave_0_readdatavalid;                                               // prio_arbiter_0:AVS_S3_READDATAVALID -> prio_arbiter_0_s3_translator:av_readdatavalid
	wire    [3:0] prio_arbiter_0_s3_translator_avalon_anti_slave_0_byteenable;                                                  // prio_arbiter_0_s3_translator:av_byteenable -> prio_arbiter_0:AVS_S3_BYTEENABLE
	wire          com_nios_instruction_master_translator_avalon_universal_master_0_waitrequest;                                 // com_nios_instruction_master_translator_avalon_universal_master_0_agent:av_waitrequest -> com_nios_instruction_master_translator:uav_waitrequest
	wire    [5:0] com_nios_instruction_master_translator_avalon_universal_master_0_burstcount;                                  // com_nios_instruction_master_translator:uav_burstcount -> com_nios_instruction_master_translator_avalon_universal_master_0_agent:av_burstcount
	wire   [31:0] com_nios_instruction_master_translator_avalon_universal_master_0_writedata;                                   // com_nios_instruction_master_translator:uav_writedata -> com_nios_instruction_master_translator_avalon_universal_master_0_agent:av_writedata
	wire   [31:0] com_nios_instruction_master_translator_avalon_universal_master_0_address;                                     // com_nios_instruction_master_translator:uav_address -> com_nios_instruction_master_translator_avalon_universal_master_0_agent:av_address
	wire          com_nios_instruction_master_translator_avalon_universal_master_0_lock;                                        // com_nios_instruction_master_translator:uav_lock -> com_nios_instruction_master_translator_avalon_universal_master_0_agent:av_lock
	wire          com_nios_instruction_master_translator_avalon_universal_master_0_write;                                       // com_nios_instruction_master_translator:uav_write -> com_nios_instruction_master_translator_avalon_universal_master_0_agent:av_write
	wire          com_nios_instruction_master_translator_avalon_universal_master_0_read;                                        // com_nios_instruction_master_translator:uav_read -> com_nios_instruction_master_translator_avalon_universal_master_0_agent:av_read
	wire   [31:0] com_nios_instruction_master_translator_avalon_universal_master_0_readdata;                                    // com_nios_instruction_master_translator_avalon_universal_master_0_agent:av_readdata -> com_nios_instruction_master_translator:uav_readdata
	wire          com_nios_instruction_master_translator_avalon_universal_master_0_debugaccess;                                 // com_nios_instruction_master_translator:uav_debugaccess -> com_nios_instruction_master_translator_avalon_universal_master_0_agent:av_debugaccess
	wire    [3:0] com_nios_instruction_master_translator_avalon_universal_master_0_byteenable;                                  // com_nios_instruction_master_translator:uav_byteenable -> com_nios_instruction_master_translator_avalon_universal_master_0_agent:av_byteenable
	wire          com_nios_instruction_master_translator_avalon_universal_master_0_readdatavalid;                               // com_nios_instruction_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> com_nios_instruction_master_translator:uav_readdatavalid
	wire          com_nios_data_master_translator_avalon_universal_master_0_waitrequest;                                        // com_nios_data_master_translator_avalon_universal_master_0_agent:av_waitrequest -> com_nios_data_master_translator:uav_waitrequest
	wire    [5:0] com_nios_data_master_translator_avalon_universal_master_0_burstcount;                                         // com_nios_data_master_translator:uav_burstcount -> com_nios_data_master_translator_avalon_universal_master_0_agent:av_burstcount
	wire   [31:0] com_nios_data_master_translator_avalon_universal_master_0_writedata;                                          // com_nios_data_master_translator:uav_writedata -> com_nios_data_master_translator_avalon_universal_master_0_agent:av_writedata
	wire   [31:0] com_nios_data_master_translator_avalon_universal_master_0_address;                                            // com_nios_data_master_translator:uav_address -> com_nios_data_master_translator_avalon_universal_master_0_agent:av_address
	wire          com_nios_data_master_translator_avalon_universal_master_0_lock;                                               // com_nios_data_master_translator:uav_lock -> com_nios_data_master_translator_avalon_universal_master_0_agent:av_lock
	wire          com_nios_data_master_translator_avalon_universal_master_0_write;                                              // com_nios_data_master_translator:uav_write -> com_nios_data_master_translator_avalon_universal_master_0_agent:av_write
	wire          com_nios_data_master_translator_avalon_universal_master_0_read;                                               // com_nios_data_master_translator:uav_read -> com_nios_data_master_translator_avalon_universal_master_0_agent:av_read
	wire   [31:0] com_nios_data_master_translator_avalon_universal_master_0_readdata;                                           // com_nios_data_master_translator_avalon_universal_master_0_agent:av_readdata -> com_nios_data_master_translator:uav_readdata
	wire          com_nios_data_master_translator_avalon_universal_master_0_debugaccess;                                        // com_nios_data_master_translator:uav_debugaccess -> com_nios_data_master_translator_avalon_universal_master_0_agent:av_debugaccess
	wire    [3:0] com_nios_data_master_translator_avalon_universal_master_0_byteenable;                                         // com_nios_data_master_translator:uav_byteenable -> com_nios_data_master_translator_avalon_universal_master_0_agent:av_byteenable
	wire          com_nios_data_master_translator_avalon_universal_master_0_readdatavalid;                                      // com_nios_data_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> com_nios_data_master_translator:uav_readdatavalid
	wire          carcontrol_nios_data_master_translator_avalon_universal_master_0_waitrequest;                                 // carControl_nios_data_master_translator_avalon_universal_master_0_agent:av_waitrequest -> carControl_nios_data_master_translator:uav_waitrequest
	wire    [2:0] carcontrol_nios_data_master_translator_avalon_universal_master_0_burstcount;                                  // carControl_nios_data_master_translator:uav_burstcount -> carControl_nios_data_master_translator_avalon_universal_master_0_agent:av_burstcount
	wire   [31:0] carcontrol_nios_data_master_translator_avalon_universal_master_0_writedata;                                   // carControl_nios_data_master_translator:uav_writedata -> carControl_nios_data_master_translator_avalon_universal_master_0_agent:av_writedata
	wire   [31:0] carcontrol_nios_data_master_translator_avalon_universal_master_0_address;                                     // carControl_nios_data_master_translator:uav_address -> carControl_nios_data_master_translator_avalon_universal_master_0_agent:av_address
	wire          carcontrol_nios_data_master_translator_avalon_universal_master_0_lock;                                        // carControl_nios_data_master_translator:uav_lock -> carControl_nios_data_master_translator_avalon_universal_master_0_agent:av_lock
	wire          carcontrol_nios_data_master_translator_avalon_universal_master_0_write;                                       // carControl_nios_data_master_translator:uav_write -> carControl_nios_data_master_translator_avalon_universal_master_0_agent:av_write
	wire          carcontrol_nios_data_master_translator_avalon_universal_master_0_read;                                        // carControl_nios_data_master_translator:uav_read -> carControl_nios_data_master_translator_avalon_universal_master_0_agent:av_read
	wire   [31:0] carcontrol_nios_data_master_translator_avalon_universal_master_0_readdata;                                    // carControl_nios_data_master_translator_avalon_universal_master_0_agent:av_readdata -> carControl_nios_data_master_translator:uav_readdata
	wire          carcontrol_nios_data_master_translator_avalon_universal_master_0_debugaccess;                                 // carControl_nios_data_master_translator:uav_debugaccess -> carControl_nios_data_master_translator_avalon_universal_master_0_agent:av_debugaccess
	wire    [3:0] carcontrol_nios_data_master_translator_avalon_universal_master_0_byteenable;                                  // carControl_nios_data_master_translator:uav_byteenable -> carControl_nios_data_master_translator_avalon_universal_master_0_agent:av_byteenable
	wire          carcontrol_nios_data_master_translator_avalon_universal_master_0_readdatavalid;                               // carControl_nios_data_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> carControl_nios_data_master_translator:uav_readdatavalid
	wire          carcontrol_nios_instruction_master_translator_avalon_universal_master_0_waitrequest;                          // carControl_nios_instruction_master_translator_avalon_universal_master_0_agent:av_waitrequest -> carControl_nios_instruction_master_translator:uav_waitrequest
	wire    [2:0] carcontrol_nios_instruction_master_translator_avalon_universal_master_0_burstcount;                           // carControl_nios_instruction_master_translator:uav_burstcount -> carControl_nios_instruction_master_translator_avalon_universal_master_0_agent:av_burstcount
	wire   [31:0] carcontrol_nios_instruction_master_translator_avalon_universal_master_0_writedata;                            // carControl_nios_instruction_master_translator:uav_writedata -> carControl_nios_instruction_master_translator_avalon_universal_master_0_agent:av_writedata
	wire   [31:0] carcontrol_nios_instruction_master_translator_avalon_universal_master_0_address;                              // carControl_nios_instruction_master_translator:uav_address -> carControl_nios_instruction_master_translator_avalon_universal_master_0_agent:av_address
	wire          carcontrol_nios_instruction_master_translator_avalon_universal_master_0_lock;                                 // carControl_nios_instruction_master_translator:uav_lock -> carControl_nios_instruction_master_translator_avalon_universal_master_0_agent:av_lock
	wire          carcontrol_nios_instruction_master_translator_avalon_universal_master_0_write;                                // carControl_nios_instruction_master_translator:uav_write -> carControl_nios_instruction_master_translator_avalon_universal_master_0_agent:av_write
	wire          carcontrol_nios_instruction_master_translator_avalon_universal_master_0_read;                                 // carControl_nios_instruction_master_translator:uav_read -> carControl_nios_instruction_master_translator_avalon_universal_master_0_agent:av_read
	wire   [31:0] carcontrol_nios_instruction_master_translator_avalon_universal_master_0_readdata;                             // carControl_nios_instruction_master_translator_avalon_universal_master_0_agent:av_readdata -> carControl_nios_instruction_master_translator:uav_readdata
	wire          carcontrol_nios_instruction_master_translator_avalon_universal_master_0_debugaccess;                          // carControl_nios_instruction_master_translator:uav_debugaccess -> carControl_nios_instruction_master_translator_avalon_universal_master_0_agent:av_debugaccess
	wire    [3:0] carcontrol_nios_instruction_master_translator_avalon_universal_master_0_byteenable;                           // carControl_nios_instruction_master_translator:uav_byteenable -> carControl_nios_instruction_master_translator_avalon_universal_master_0_agent:av_byteenable
	wire          carcontrol_nios_instruction_master_translator_avalon_universal_master_0_readdatavalid;                        // carControl_nios_instruction_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> carControl_nios_instruction_master_translator:uav_readdatavalid
	wire          ethernet_subsystem_sgdma_rx_m_write_translator_avalon_universal_master_0_waitrequest;                         // ethernet_subsystem_sgdma_rx_m_write_translator_avalon_universal_master_0_agent:av_waitrequest -> ethernet_subsystem_sgdma_rx_m_write_translator:uav_waitrequest
	wire    [2:0] ethernet_subsystem_sgdma_rx_m_write_translator_avalon_universal_master_0_burstcount;                          // ethernet_subsystem_sgdma_rx_m_write_translator:uav_burstcount -> ethernet_subsystem_sgdma_rx_m_write_translator_avalon_universal_master_0_agent:av_burstcount
	wire   [31:0] ethernet_subsystem_sgdma_rx_m_write_translator_avalon_universal_master_0_writedata;                           // ethernet_subsystem_sgdma_rx_m_write_translator:uav_writedata -> ethernet_subsystem_sgdma_rx_m_write_translator_avalon_universal_master_0_agent:av_writedata
	wire   [31:0] ethernet_subsystem_sgdma_rx_m_write_translator_avalon_universal_master_0_address;                             // ethernet_subsystem_sgdma_rx_m_write_translator:uav_address -> ethernet_subsystem_sgdma_rx_m_write_translator_avalon_universal_master_0_agent:av_address
	wire          ethernet_subsystem_sgdma_rx_m_write_translator_avalon_universal_master_0_lock;                                // ethernet_subsystem_sgdma_rx_m_write_translator:uav_lock -> ethernet_subsystem_sgdma_rx_m_write_translator_avalon_universal_master_0_agent:av_lock
	wire          ethernet_subsystem_sgdma_rx_m_write_translator_avalon_universal_master_0_write;                               // ethernet_subsystem_sgdma_rx_m_write_translator:uav_write -> ethernet_subsystem_sgdma_rx_m_write_translator_avalon_universal_master_0_agent:av_write
	wire          ethernet_subsystem_sgdma_rx_m_write_translator_avalon_universal_master_0_read;                                // ethernet_subsystem_sgdma_rx_m_write_translator:uav_read -> ethernet_subsystem_sgdma_rx_m_write_translator_avalon_universal_master_0_agent:av_read
	wire   [31:0] ethernet_subsystem_sgdma_rx_m_write_translator_avalon_universal_master_0_readdata;                            // ethernet_subsystem_sgdma_rx_m_write_translator_avalon_universal_master_0_agent:av_readdata -> ethernet_subsystem_sgdma_rx_m_write_translator:uav_readdata
	wire          ethernet_subsystem_sgdma_rx_m_write_translator_avalon_universal_master_0_debugaccess;                         // ethernet_subsystem_sgdma_rx_m_write_translator:uav_debugaccess -> ethernet_subsystem_sgdma_rx_m_write_translator_avalon_universal_master_0_agent:av_debugaccess
	wire    [3:0] ethernet_subsystem_sgdma_rx_m_write_translator_avalon_universal_master_0_byteenable;                          // ethernet_subsystem_sgdma_rx_m_write_translator:uav_byteenable -> ethernet_subsystem_sgdma_rx_m_write_translator_avalon_universal_master_0_agent:av_byteenable
	wire          ethernet_subsystem_sgdma_rx_m_write_translator_avalon_universal_master_0_readdatavalid;                       // ethernet_subsystem_sgdma_rx_m_write_translator_avalon_universal_master_0_agent:av_readdatavalid -> ethernet_subsystem_sgdma_rx_m_write_translator:uav_readdatavalid
	wire          ethernet_subsystem_sgdma_tx_m_read_translator_avalon_universal_master_0_waitrequest;                          // ethernet_subsystem_sgdma_tx_m_read_translator_avalon_universal_master_0_agent:av_waitrequest -> ethernet_subsystem_sgdma_tx_m_read_translator:uav_waitrequest
	wire    [2:0] ethernet_subsystem_sgdma_tx_m_read_translator_avalon_universal_master_0_burstcount;                           // ethernet_subsystem_sgdma_tx_m_read_translator:uav_burstcount -> ethernet_subsystem_sgdma_tx_m_read_translator_avalon_universal_master_0_agent:av_burstcount
	wire   [31:0] ethernet_subsystem_sgdma_tx_m_read_translator_avalon_universal_master_0_writedata;                            // ethernet_subsystem_sgdma_tx_m_read_translator:uav_writedata -> ethernet_subsystem_sgdma_tx_m_read_translator_avalon_universal_master_0_agent:av_writedata
	wire   [31:0] ethernet_subsystem_sgdma_tx_m_read_translator_avalon_universal_master_0_address;                              // ethernet_subsystem_sgdma_tx_m_read_translator:uav_address -> ethernet_subsystem_sgdma_tx_m_read_translator_avalon_universal_master_0_agent:av_address
	wire          ethernet_subsystem_sgdma_tx_m_read_translator_avalon_universal_master_0_lock;                                 // ethernet_subsystem_sgdma_tx_m_read_translator:uav_lock -> ethernet_subsystem_sgdma_tx_m_read_translator_avalon_universal_master_0_agent:av_lock
	wire          ethernet_subsystem_sgdma_tx_m_read_translator_avalon_universal_master_0_write;                                // ethernet_subsystem_sgdma_tx_m_read_translator:uav_write -> ethernet_subsystem_sgdma_tx_m_read_translator_avalon_universal_master_0_agent:av_write
	wire          ethernet_subsystem_sgdma_tx_m_read_translator_avalon_universal_master_0_read;                                 // ethernet_subsystem_sgdma_tx_m_read_translator:uav_read -> ethernet_subsystem_sgdma_tx_m_read_translator_avalon_universal_master_0_agent:av_read
	wire   [31:0] ethernet_subsystem_sgdma_tx_m_read_translator_avalon_universal_master_0_readdata;                             // ethernet_subsystem_sgdma_tx_m_read_translator_avalon_universal_master_0_agent:av_readdata -> ethernet_subsystem_sgdma_tx_m_read_translator:uav_readdata
	wire          ethernet_subsystem_sgdma_tx_m_read_translator_avalon_universal_master_0_debugaccess;                          // ethernet_subsystem_sgdma_tx_m_read_translator:uav_debugaccess -> ethernet_subsystem_sgdma_tx_m_read_translator_avalon_universal_master_0_agent:av_debugaccess
	wire    [3:0] ethernet_subsystem_sgdma_tx_m_read_translator_avalon_universal_master_0_byteenable;                           // ethernet_subsystem_sgdma_tx_m_read_translator:uav_byteenable -> ethernet_subsystem_sgdma_tx_m_read_translator_avalon_universal_master_0_agent:av_byteenable
	wire          ethernet_subsystem_sgdma_tx_m_read_translator_avalon_universal_master_0_readdatavalid;                        // ethernet_subsystem_sgdma_tx_m_read_translator_avalon_universal_master_0_agent:av_readdatavalid -> ethernet_subsystem_sgdma_tx_m_read_translator:uav_readdatavalid
	wire          com_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest;                          // com_nios_jtag_debug_module_translator:uav_waitrequest -> com_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] com_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount;                           // com_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_burstcount -> com_nios_jtag_debug_module_translator:uav_burstcount
	wire   [31:0] com_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata;                            // com_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_writedata -> com_nios_jtag_debug_module_translator:uav_writedata
	wire   [31:0] com_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address;                              // com_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_address -> com_nios_jtag_debug_module_translator:uav_address
	wire          com_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write;                                // com_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_write -> com_nios_jtag_debug_module_translator:uav_write
	wire          com_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock;                                 // com_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_lock -> com_nios_jtag_debug_module_translator:uav_lock
	wire          com_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read;                                 // com_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_read -> com_nios_jtag_debug_module_translator:uav_read
	wire   [31:0] com_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata;                             // com_nios_jtag_debug_module_translator:uav_readdata -> com_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          com_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                        // com_nios_jtag_debug_module_translator:uav_readdatavalid -> com_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          com_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess;                          // com_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_debugaccess -> com_nios_jtag_debug_module_translator:uav_debugaccess
	wire    [3:0] com_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable;                           // com_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_byteenable -> com_nios_jtag_debug_module_translator:uav_byteenable
	wire          com_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                   // com_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> com_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          com_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid;                         // com_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_valid -> com_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          com_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                 // com_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> com_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [113:0] com_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data;                          // com_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_data -> com_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          com_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready;                         // com_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> com_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          com_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                // com_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> com_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          com_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                      // com_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> com_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          com_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;              // com_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> com_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [113:0] com_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                       // com_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> com_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          com_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                      // com_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_ready -> com_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          com_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                    // com_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> com_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] com_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                     // com_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> com_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          com_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                    // com_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> com_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          com_memory_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                       // com_memory_s1_translator:uav_waitrequest -> com_memory_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] com_memory_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                        // com_memory_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> com_memory_s1_translator:uav_burstcount
	wire   [31:0] com_memory_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                         // com_memory_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> com_memory_s1_translator:uav_writedata
	wire   [31:0] com_memory_s1_translator_avalon_universal_slave_0_agent_m0_address;                                           // com_memory_s1_translator_avalon_universal_slave_0_agent:m0_address -> com_memory_s1_translator:uav_address
	wire          com_memory_s1_translator_avalon_universal_slave_0_agent_m0_write;                                             // com_memory_s1_translator_avalon_universal_slave_0_agent:m0_write -> com_memory_s1_translator:uav_write
	wire          com_memory_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                              // com_memory_s1_translator_avalon_universal_slave_0_agent:m0_lock -> com_memory_s1_translator:uav_lock
	wire          com_memory_s1_translator_avalon_universal_slave_0_agent_m0_read;                                              // com_memory_s1_translator_avalon_universal_slave_0_agent:m0_read -> com_memory_s1_translator:uav_read
	wire   [31:0] com_memory_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                          // com_memory_s1_translator:uav_readdata -> com_memory_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          com_memory_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                     // com_memory_s1_translator:uav_readdatavalid -> com_memory_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          com_memory_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                       // com_memory_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> com_memory_s1_translator:uav_debugaccess
	wire    [3:0] com_memory_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                        // com_memory_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> com_memory_s1_translator:uav_byteenable
	wire          com_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                                // com_memory_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> com_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          com_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                      // com_memory_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> com_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          com_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                              // com_memory_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> com_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [113:0] com_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                       // com_memory_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> com_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          com_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                      // com_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> com_memory_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          com_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                             // com_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> com_memory_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          com_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                   // com_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> com_memory_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          com_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                           // com_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> com_memory_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [113:0] com_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                    // com_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> com_memory_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          com_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                   // com_memory_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> com_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          com_memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                                 // com_memory_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> com_memory_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] com_memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                                  // com_memory_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> com_memory_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          com_memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                                 // com_memory_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> com_memory_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          jtaguart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;                        // jtaguart_0_avalon_jtag_slave_translator:uav_waitrequest -> jtaguart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] jtaguart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;                         // jtaguart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> jtaguart_0_avalon_jtag_slave_translator:uav_burstcount
	wire   [31:0] jtaguart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata;                          // jtaguart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> jtaguart_0_avalon_jtag_slave_translator:uav_writedata
	wire   [31:0] jtaguart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address;                            // jtaguart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_address -> jtaguart_0_avalon_jtag_slave_translator:uav_address
	wire          jtaguart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write;                              // jtaguart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_write -> jtaguart_0_avalon_jtag_slave_translator:uav_write
	wire          jtaguart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock;                               // jtaguart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_lock -> jtaguart_0_avalon_jtag_slave_translator:uav_lock
	wire          jtaguart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read;                               // jtaguart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_read -> jtaguart_0_avalon_jtag_slave_translator:uav_read
	wire   [31:0] jtaguart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                           // jtaguart_0_avalon_jtag_slave_translator:uav_readdata -> jtaguart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          jtaguart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                      // jtaguart_0_avalon_jtag_slave_translator:uav_readdatavalid -> jtaguart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          jtaguart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;                        // jtaguart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> jtaguart_0_avalon_jtag_slave_translator:uav_debugaccess
	wire    [3:0] jtaguart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;                         // jtaguart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> jtaguart_0_avalon_jtag_slave_translator:uav_byteenable
	wire          jtaguart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                 // jtaguart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> jtaguart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          jtaguart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;                       // jtaguart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> jtaguart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          jtaguart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;               // jtaguart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> jtaguart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [113:0] jtaguart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data;                        // jtaguart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> jtaguart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          jtaguart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;                       // jtaguart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> jtaguart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          jtaguart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;              // jtaguart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> jtaguart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          jtaguart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                    // jtaguart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> jtaguart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          jtaguart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;            // jtaguart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> jtaguart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [113:0] jtaguart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                     // jtaguart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> jtaguart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          jtaguart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                    // jtaguart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> jtaguart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          jtaguart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                  // jtaguart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> jtaguart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] jtaguart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                   // jtaguart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> jtaguart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          jtaguart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                  // jtaguart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> jtaguart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          shared_memory_mutex_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                              // shared_memory_mutex_s1_translator:uav_waitrequest -> shared_memory_mutex_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] shared_memory_mutex_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                               // shared_memory_mutex_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> shared_memory_mutex_s1_translator:uav_burstcount
	wire   [31:0] shared_memory_mutex_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                // shared_memory_mutex_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> shared_memory_mutex_s1_translator:uav_writedata
	wire   [31:0] shared_memory_mutex_s1_translator_avalon_universal_slave_0_agent_m0_address;                                  // shared_memory_mutex_s1_translator_avalon_universal_slave_0_agent:m0_address -> shared_memory_mutex_s1_translator:uav_address
	wire          shared_memory_mutex_s1_translator_avalon_universal_slave_0_agent_m0_write;                                    // shared_memory_mutex_s1_translator_avalon_universal_slave_0_agent:m0_write -> shared_memory_mutex_s1_translator:uav_write
	wire          shared_memory_mutex_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                     // shared_memory_mutex_s1_translator_avalon_universal_slave_0_agent:m0_lock -> shared_memory_mutex_s1_translator:uav_lock
	wire          shared_memory_mutex_s1_translator_avalon_universal_slave_0_agent_m0_read;                                     // shared_memory_mutex_s1_translator_avalon_universal_slave_0_agent:m0_read -> shared_memory_mutex_s1_translator:uav_read
	wire   [31:0] shared_memory_mutex_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                 // shared_memory_mutex_s1_translator:uav_readdata -> shared_memory_mutex_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          shared_memory_mutex_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                            // shared_memory_mutex_s1_translator:uav_readdatavalid -> shared_memory_mutex_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          shared_memory_mutex_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                              // shared_memory_mutex_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> shared_memory_mutex_s1_translator:uav_debugaccess
	wire    [3:0] shared_memory_mutex_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                               // shared_memory_mutex_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> shared_memory_mutex_s1_translator:uav_byteenable
	wire          shared_memory_mutex_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                       // shared_memory_mutex_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> shared_memory_mutex_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          shared_memory_mutex_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                             // shared_memory_mutex_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> shared_memory_mutex_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          shared_memory_mutex_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                     // shared_memory_mutex_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> shared_memory_mutex_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [113:0] shared_memory_mutex_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                              // shared_memory_mutex_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> shared_memory_mutex_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          shared_memory_mutex_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                             // shared_memory_mutex_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> shared_memory_mutex_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          shared_memory_mutex_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                    // shared_memory_mutex_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> shared_memory_mutex_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          shared_memory_mutex_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                          // shared_memory_mutex_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> shared_memory_mutex_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          shared_memory_mutex_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                  // shared_memory_mutex_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> shared_memory_mutex_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [113:0] shared_memory_mutex_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                           // shared_memory_mutex_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> shared_memory_mutex_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          shared_memory_mutex_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                          // shared_memory_mutex_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> shared_memory_mutex_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          shared_memory_mutex_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                        // shared_memory_mutex_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> shared_memory_mutex_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] shared_memory_mutex_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                         // shared_memory_mutex_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> shared_memory_mutex_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          shared_memory_mutex_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                        // shared_memory_mutex_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> shared_memory_mutex_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          com_timer_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                        // com_timer_s1_translator:uav_waitrequest -> com_timer_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] com_timer_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                         // com_timer_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> com_timer_s1_translator:uav_burstcount
	wire   [31:0] com_timer_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                          // com_timer_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> com_timer_s1_translator:uav_writedata
	wire   [31:0] com_timer_s1_translator_avalon_universal_slave_0_agent_m0_address;                                            // com_timer_s1_translator_avalon_universal_slave_0_agent:m0_address -> com_timer_s1_translator:uav_address
	wire          com_timer_s1_translator_avalon_universal_slave_0_agent_m0_write;                                              // com_timer_s1_translator_avalon_universal_slave_0_agent:m0_write -> com_timer_s1_translator:uav_write
	wire          com_timer_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                               // com_timer_s1_translator_avalon_universal_slave_0_agent:m0_lock -> com_timer_s1_translator:uav_lock
	wire          com_timer_s1_translator_avalon_universal_slave_0_agent_m0_read;                                               // com_timer_s1_translator_avalon_universal_slave_0_agent:m0_read -> com_timer_s1_translator:uav_read
	wire   [31:0] com_timer_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                           // com_timer_s1_translator:uav_readdata -> com_timer_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          com_timer_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                      // com_timer_s1_translator:uav_readdatavalid -> com_timer_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          com_timer_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                        // com_timer_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> com_timer_s1_translator:uav_debugaccess
	wire    [3:0] com_timer_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                         // com_timer_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> com_timer_s1_translator:uav_byteenable
	wire          com_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                                 // com_timer_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> com_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          com_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                       // com_timer_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> com_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          com_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                               // com_timer_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> com_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [113:0] com_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                        // com_timer_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> com_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          com_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                       // com_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> com_timer_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          com_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                              // com_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> com_timer_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          com_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                    // com_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> com_timer_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          com_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                            // com_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> com_timer_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [113:0] com_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                     // com_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> com_timer_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          com_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                    // com_timer_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> com_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          com_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                                  // com_timer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> com_timer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] com_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                                   // com_timer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> com_timer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          com_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                                  // com_timer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> com_timer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          ethernet_subsystem_ethernet_bridge_s0_translator_avalon_universal_slave_0_agent_m0_waitrequest;               // ethernet_subsystem_ethernet_bridge_s0_translator:uav_waitrequest -> ethernet_subsystem_ethernet_bridge_s0_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] ethernet_subsystem_ethernet_bridge_s0_translator_avalon_universal_slave_0_agent_m0_burstcount;                // ethernet_subsystem_ethernet_bridge_s0_translator_avalon_universal_slave_0_agent:m0_burstcount -> ethernet_subsystem_ethernet_bridge_s0_translator:uav_burstcount
	wire   [31:0] ethernet_subsystem_ethernet_bridge_s0_translator_avalon_universal_slave_0_agent_m0_writedata;                 // ethernet_subsystem_ethernet_bridge_s0_translator_avalon_universal_slave_0_agent:m0_writedata -> ethernet_subsystem_ethernet_bridge_s0_translator:uav_writedata
	wire   [31:0] ethernet_subsystem_ethernet_bridge_s0_translator_avalon_universal_slave_0_agent_m0_address;                   // ethernet_subsystem_ethernet_bridge_s0_translator_avalon_universal_slave_0_agent:m0_address -> ethernet_subsystem_ethernet_bridge_s0_translator:uav_address
	wire          ethernet_subsystem_ethernet_bridge_s0_translator_avalon_universal_slave_0_agent_m0_write;                     // ethernet_subsystem_ethernet_bridge_s0_translator_avalon_universal_slave_0_agent:m0_write -> ethernet_subsystem_ethernet_bridge_s0_translator:uav_write
	wire          ethernet_subsystem_ethernet_bridge_s0_translator_avalon_universal_slave_0_agent_m0_lock;                      // ethernet_subsystem_ethernet_bridge_s0_translator_avalon_universal_slave_0_agent:m0_lock -> ethernet_subsystem_ethernet_bridge_s0_translator:uav_lock
	wire          ethernet_subsystem_ethernet_bridge_s0_translator_avalon_universal_slave_0_agent_m0_read;                      // ethernet_subsystem_ethernet_bridge_s0_translator_avalon_universal_slave_0_agent:m0_read -> ethernet_subsystem_ethernet_bridge_s0_translator:uav_read
	wire   [31:0] ethernet_subsystem_ethernet_bridge_s0_translator_avalon_universal_slave_0_agent_m0_readdata;                  // ethernet_subsystem_ethernet_bridge_s0_translator:uav_readdata -> ethernet_subsystem_ethernet_bridge_s0_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          ethernet_subsystem_ethernet_bridge_s0_translator_avalon_universal_slave_0_agent_m0_readdatavalid;             // ethernet_subsystem_ethernet_bridge_s0_translator:uav_readdatavalid -> ethernet_subsystem_ethernet_bridge_s0_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          ethernet_subsystem_ethernet_bridge_s0_translator_avalon_universal_slave_0_agent_m0_debugaccess;               // ethernet_subsystem_ethernet_bridge_s0_translator_avalon_universal_slave_0_agent:m0_debugaccess -> ethernet_subsystem_ethernet_bridge_s0_translator:uav_debugaccess
	wire    [3:0] ethernet_subsystem_ethernet_bridge_s0_translator_avalon_universal_slave_0_agent_m0_byteenable;                // ethernet_subsystem_ethernet_bridge_s0_translator_avalon_universal_slave_0_agent:m0_byteenable -> ethernet_subsystem_ethernet_bridge_s0_translator:uav_byteenable
	wire          ethernet_subsystem_ethernet_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;        // ethernet_subsystem_ethernet_bridge_s0_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> ethernet_subsystem_ethernet_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          ethernet_subsystem_ethernet_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_valid;              // ethernet_subsystem_ethernet_bridge_s0_translator_avalon_universal_slave_0_agent:rf_source_valid -> ethernet_subsystem_ethernet_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          ethernet_subsystem_ethernet_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;      // ethernet_subsystem_ethernet_bridge_s0_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> ethernet_subsystem_ethernet_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [113:0] ethernet_subsystem_ethernet_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_data;               // ethernet_subsystem_ethernet_bridge_s0_translator_avalon_universal_slave_0_agent:rf_source_data -> ethernet_subsystem_ethernet_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          ethernet_subsystem_ethernet_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_ready;              // ethernet_subsystem_ethernet_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> ethernet_subsystem_ethernet_bridge_s0_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          ethernet_subsystem_ethernet_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;     // ethernet_subsystem_ethernet_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> ethernet_subsystem_ethernet_bridge_s0_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          ethernet_subsystem_ethernet_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;           // ethernet_subsystem_ethernet_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> ethernet_subsystem_ethernet_bridge_s0_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          ethernet_subsystem_ethernet_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;   // ethernet_subsystem_ethernet_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> ethernet_subsystem_ethernet_bridge_s0_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [113:0] ethernet_subsystem_ethernet_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;            // ethernet_subsystem_ethernet_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> ethernet_subsystem_ethernet_bridge_s0_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          ethernet_subsystem_ethernet_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;           // ethernet_subsystem_ethernet_bridge_s0_translator_avalon_universal_slave_0_agent:rf_sink_ready -> ethernet_subsystem_ethernet_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          ethernet_subsystem_ethernet_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;         // ethernet_subsystem_ethernet_bridge_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> ethernet_subsystem_ethernet_bridge_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] ethernet_subsystem_ethernet_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;          // ethernet_subsystem_ethernet_bridge_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> ethernet_subsystem_ethernet_bridge_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          ethernet_subsystem_ethernet_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;         // ethernet_subsystem_ethernet_bridge_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> ethernet_subsystem_ethernet_bridge_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          ethernet_subsystem_descriptor_memory_s2_translator_avalon_universal_slave_0_agent_m0_waitrequest;             // ethernet_subsystem_descriptor_memory_s2_translator:uav_waitrequest -> ethernet_subsystem_descriptor_memory_s2_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] ethernet_subsystem_descriptor_memory_s2_translator_avalon_universal_slave_0_agent_m0_burstcount;              // ethernet_subsystem_descriptor_memory_s2_translator_avalon_universal_slave_0_agent:m0_burstcount -> ethernet_subsystem_descriptor_memory_s2_translator:uav_burstcount
	wire   [31:0] ethernet_subsystem_descriptor_memory_s2_translator_avalon_universal_slave_0_agent_m0_writedata;               // ethernet_subsystem_descriptor_memory_s2_translator_avalon_universal_slave_0_agent:m0_writedata -> ethernet_subsystem_descriptor_memory_s2_translator:uav_writedata
	wire   [31:0] ethernet_subsystem_descriptor_memory_s2_translator_avalon_universal_slave_0_agent_m0_address;                 // ethernet_subsystem_descriptor_memory_s2_translator_avalon_universal_slave_0_agent:m0_address -> ethernet_subsystem_descriptor_memory_s2_translator:uav_address
	wire          ethernet_subsystem_descriptor_memory_s2_translator_avalon_universal_slave_0_agent_m0_write;                   // ethernet_subsystem_descriptor_memory_s2_translator_avalon_universal_slave_0_agent:m0_write -> ethernet_subsystem_descriptor_memory_s2_translator:uav_write
	wire          ethernet_subsystem_descriptor_memory_s2_translator_avalon_universal_slave_0_agent_m0_lock;                    // ethernet_subsystem_descriptor_memory_s2_translator_avalon_universal_slave_0_agent:m0_lock -> ethernet_subsystem_descriptor_memory_s2_translator:uav_lock
	wire          ethernet_subsystem_descriptor_memory_s2_translator_avalon_universal_slave_0_agent_m0_read;                    // ethernet_subsystem_descriptor_memory_s2_translator_avalon_universal_slave_0_agent:m0_read -> ethernet_subsystem_descriptor_memory_s2_translator:uav_read
	wire   [31:0] ethernet_subsystem_descriptor_memory_s2_translator_avalon_universal_slave_0_agent_m0_readdata;                // ethernet_subsystem_descriptor_memory_s2_translator:uav_readdata -> ethernet_subsystem_descriptor_memory_s2_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          ethernet_subsystem_descriptor_memory_s2_translator_avalon_universal_slave_0_agent_m0_readdatavalid;           // ethernet_subsystem_descriptor_memory_s2_translator:uav_readdatavalid -> ethernet_subsystem_descriptor_memory_s2_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          ethernet_subsystem_descriptor_memory_s2_translator_avalon_universal_slave_0_agent_m0_debugaccess;             // ethernet_subsystem_descriptor_memory_s2_translator_avalon_universal_slave_0_agent:m0_debugaccess -> ethernet_subsystem_descriptor_memory_s2_translator:uav_debugaccess
	wire    [3:0] ethernet_subsystem_descriptor_memory_s2_translator_avalon_universal_slave_0_agent_m0_byteenable;              // ethernet_subsystem_descriptor_memory_s2_translator_avalon_universal_slave_0_agent:m0_byteenable -> ethernet_subsystem_descriptor_memory_s2_translator:uav_byteenable
	wire          ethernet_subsystem_descriptor_memory_s2_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;      // ethernet_subsystem_descriptor_memory_s2_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> ethernet_subsystem_descriptor_memory_s2_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          ethernet_subsystem_descriptor_memory_s2_translator_avalon_universal_slave_0_agent_rf_source_valid;            // ethernet_subsystem_descriptor_memory_s2_translator_avalon_universal_slave_0_agent:rf_source_valid -> ethernet_subsystem_descriptor_memory_s2_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          ethernet_subsystem_descriptor_memory_s2_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;    // ethernet_subsystem_descriptor_memory_s2_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> ethernet_subsystem_descriptor_memory_s2_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [113:0] ethernet_subsystem_descriptor_memory_s2_translator_avalon_universal_slave_0_agent_rf_source_data;             // ethernet_subsystem_descriptor_memory_s2_translator_avalon_universal_slave_0_agent:rf_source_data -> ethernet_subsystem_descriptor_memory_s2_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          ethernet_subsystem_descriptor_memory_s2_translator_avalon_universal_slave_0_agent_rf_source_ready;            // ethernet_subsystem_descriptor_memory_s2_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> ethernet_subsystem_descriptor_memory_s2_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          ethernet_subsystem_descriptor_memory_s2_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;   // ethernet_subsystem_descriptor_memory_s2_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> ethernet_subsystem_descriptor_memory_s2_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          ethernet_subsystem_descriptor_memory_s2_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;         // ethernet_subsystem_descriptor_memory_s2_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> ethernet_subsystem_descriptor_memory_s2_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          ethernet_subsystem_descriptor_memory_s2_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket; // ethernet_subsystem_descriptor_memory_s2_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> ethernet_subsystem_descriptor_memory_s2_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [113:0] ethernet_subsystem_descriptor_memory_s2_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;          // ethernet_subsystem_descriptor_memory_s2_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> ethernet_subsystem_descriptor_memory_s2_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          ethernet_subsystem_descriptor_memory_s2_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;         // ethernet_subsystem_descriptor_memory_s2_translator_avalon_universal_slave_0_agent:rf_sink_ready -> ethernet_subsystem_descriptor_memory_s2_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          ethernet_subsystem_descriptor_memory_s2_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;       // ethernet_subsystem_descriptor_memory_s2_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> ethernet_subsystem_descriptor_memory_s2_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] ethernet_subsystem_descriptor_memory_s2_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;        // ethernet_subsystem_descriptor_memory_s2_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> ethernet_subsystem_descriptor_memory_s2_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          ethernet_subsystem_descriptor_memory_s2_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;       // ethernet_subsystem_descriptor_memory_s2_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> ethernet_subsystem_descriptor_memory_s2_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          prio_arbiter_0_s0_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                   // prio_arbiter_0_s0_translator:uav_waitrequest -> prio_arbiter_0_s0_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] prio_arbiter_0_s0_translator_avalon_universal_slave_0_agent_m0_burstcount;                                    // prio_arbiter_0_s0_translator_avalon_universal_slave_0_agent:m0_burstcount -> prio_arbiter_0_s0_translator:uav_burstcount
	wire   [31:0] prio_arbiter_0_s0_translator_avalon_universal_slave_0_agent_m0_writedata;                                     // prio_arbiter_0_s0_translator_avalon_universal_slave_0_agent:m0_writedata -> prio_arbiter_0_s0_translator:uav_writedata
	wire   [31:0] prio_arbiter_0_s0_translator_avalon_universal_slave_0_agent_m0_address;                                       // prio_arbiter_0_s0_translator_avalon_universal_slave_0_agent:m0_address -> prio_arbiter_0_s0_translator:uav_address
	wire          prio_arbiter_0_s0_translator_avalon_universal_slave_0_agent_m0_write;                                         // prio_arbiter_0_s0_translator_avalon_universal_slave_0_agent:m0_write -> prio_arbiter_0_s0_translator:uav_write
	wire          prio_arbiter_0_s0_translator_avalon_universal_slave_0_agent_m0_lock;                                          // prio_arbiter_0_s0_translator_avalon_universal_slave_0_agent:m0_lock -> prio_arbiter_0_s0_translator:uav_lock
	wire          prio_arbiter_0_s0_translator_avalon_universal_slave_0_agent_m0_read;                                          // prio_arbiter_0_s0_translator_avalon_universal_slave_0_agent:m0_read -> prio_arbiter_0_s0_translator:uav_read
	wire   [31:0] prio_arbiter_0_s0_translator_avalon_universal_slave_0_agent_m0_readdata;                                      // prio_arbiter_0_s0_translator:uav_readdata -> prio_arbiter_0_s0_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          prio_arbiter_0_s0_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                 // prio_arbiter_0_s0_translator:uav_readdatavalid -> prio_arbiter_0_s0_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          prio_arbiter_0_s0_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                   // prio_arbiter_0_s0_translator_avalon_universal_slave_0_agent:m0_debugaccess -> prio_arbiter_0_s0_translator:uav_debugaccess
	wire    [3:0] prio_arbiter_0_s0_translator_avalon_universal_slave_0_agent_m0_byteenable;                                    // prio_arbiter_0_s0_translator_avalon_universal_slave_0_agent:m0_byteenable -> prio_arbiter_0_s0_translator:uav_byteenable
	wire          prio_arbiter_0_s0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                            // prio_arbiter_0_s0_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> prio_arbiter_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          prio_arbiter_0_s0_translator_avalon_universal_slave_0_agent_rf_source_valid;                                  // prio_arbiter_0_s0_translator_avalon_universal_slave_0_agent:rf_source_valid -> prio_arbiter_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          prio_arbiter_0_s0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                          // prio_arbiter_0_s0_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> prio_arbiter_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [113:0] prio_arbiter_0_s0_translator_avalon_universal_slave_0_agent_rf_source_data;                                   // prio_arbiter_0_s0_translator_avalon_universal_slave_0_agent:rf_source_data -> prio_arbiter_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          prio_arbiter_0_s0_translator_avalon_universal_slave_0_agent_rf_source_ready;                                  // prio_arbiter_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> prio_arbiter_0_s0_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          prio_arbiter_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                         // prio_arbiter_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> prio_arbiter_0_s0_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          prio_arbiter_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                               // prio_arbiter_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> prio_arbiter_0_s0_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          prio_arbiter_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                       // prio_arbiter_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> prio_arbiter_0_s0_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [113:0] prio_arbiter_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                // prio_arbiter_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> prio_arbiter_0_s0_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          prio_arbiter_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                               // prio_arbiter_0_s0_translator_avalon_universal_slave_0_agent:rf_sink_ready -> prio_arbiter_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          prio_arbiter_0_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                             // prio_arbiter_0_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> prio_arbiter_0_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] prio_arbiter_0_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                              // prio_arbiter_0_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> prio_arbiter_0_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          prio_arbiter_0_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                             // prio_arbiter_0_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> prio_arbiter_0_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          carcontrol_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest;                   // carControl_nios_jtag_debug_module_translator:uav_waitrequest -> carControl_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] carcontrol_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount;                    // carControl_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_burstcount -> carControl_nios_jtag_debug_module_translator:uav_burstcount
	wire   [31:0] carcontrol_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata;                     // carControl_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_writedata -> carControl_nios_jtag_debug_module_translator:uav_writedata
	wire   [31:0] carcontrol_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address;                       // carControl_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_address -> carControl_nios_jtag_debug_module_translator:uav_address
	wire          carcontrol_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write;                         // carControl_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_write -> carControl_nios_jtag_debug_module_translator:uav_write
	wire          carcontrol_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock;                          // carControl_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_lock -> carControl_nios_jtag_debug_module_translator:uav_lock
	wire          carcontrol_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read;                          // carControl_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_read -> carControl_nios_jtag_debug_module_translator:uav_read
	wire   [31:0] carcontrol_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata;                      // carControl_nios_jtag_debug_module_translator:uav_readdata -> carControl_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          carcontrol_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                 // carControl_nios_jtag_debug_module_translator:uav_readdatavalid -> carControl_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          carcontrol_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess;                   // carControl_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_debugaccess -> carControl_nios_jtag_debug_module_translator:uav_debugaccess
	wire    [3:0] carcontrol_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable;                    // carControl_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_byteenable -> carControl_nios_jtag_debug_module_translator:uav_byteenable
	wire          carcontrol_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;            // carControl_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> carControl_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          carcontrol_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid;                  // carControl_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_valid -> carControl_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          carcontrol_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;          // carControl_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> carControl_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [113:0] carcontrol_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data;                   // carControl_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_data -> carControl_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          carcontrol_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready;                  // carControl_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> carControl_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          carcontrol_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;         // carControl_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> carControl_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          carcontrol_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;               // carControl_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> carControl_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          carcontrol_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;       // carControl_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> carControl_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [113:0] carcontrol_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                // carControl_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> carControl_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          carcontrol_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;               // carControl_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_ready -> carControl_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          carcontrol_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;             // carControl_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> carControl_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] carcontrol_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;              // carControl_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> carControl_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          carcontrol_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;             // carControl_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> carControl_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                 // onchip_memory2_0_s1_translator:uav_waitrequest -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                  // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> onchip_memory2_0_s1_translator:uav_burstcount
	wire   [31:0] onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                   // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> onchip_memory2_0_s1_translator:uav_writedata
	wire   [31:0] onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_address;                                     // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:m0_address -> onchip_memory2_0_s1_translator:uav_address
	wire          onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_write;                                       // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:m0_write -> onchip_memory2_0_s1_translator:uav_write
	wire          onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                        // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:m0_lock -> onchip_memory2_0_s1_translator:uav_lock
	wire          onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_read;                                        // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:m0_read -> onchip_memory2_0_s1_translator:uav_read
	wire   [31:0] onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                    // onchip_memory2_0_s1_translator:uav_readdata -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                               // onchip_memory2_0_s1_translator:uav_readdatavalid -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                 // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> onchip_memory2_0_s1_translator:uav_debugaccess
	wire    [3:0] onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                  // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> onchip_memory2_0_s1_translator:uav_byteenable
	wire          onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                          // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                        // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [113:0] onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                 // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                       // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                             // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                     // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [113:0] onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                              // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                             // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                           // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                            // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                           // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          jtaguart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;                        // jtaguart_1_avalon_jtag_slave_translator:uav_waitrequest -> jtaguart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] jtaguart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;                         // jtaguart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> jtaguart_1_avalon_jtag_slave_translator:uav_burstcount
	wire   [31:0] jtaguart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata;                          // jtaguart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> jtaguart_1_avalon_jtag_slave_translator:uav_writedata
	wire   [31:0] jtaguart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address;                            // jtaguart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_address -> jtaguart_1_avalon_jtag_slave_translator:uav_address
	wire          jtaguart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write;                              // jtaguart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_write -> jtaguart_1_avalon_jtag_slave_translator:uav_write
	wire          jtaguart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock;                               // jtaguart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_lock -> jtaguart_1_avalon_jtag_slave_translator:uav_lock
	wire          jtaguart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read;                               // jtaguart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_read -> jtaguart_1_avalon_jtag_slave_translator:uav_read
	wire   [31:0] jtaguart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                           // jtaguart_1_avalon_jtag_slave_translator:uav_readdata -> jtaguart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          jtaguart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                      // jtaguart_1_avalon_jtag_slave_translator:uav_readdatavalid -> jtaguart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          jtaguart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;                        // jtaguart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> jtaguart_1_avalon_jtag_slave_translator:uav_debugaccess
	wire    [3:0] jtaguart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;                         // jtaguart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> jtaguart_1_avalon_jtag_slave_translator:uav_byteenable
	wire          jtaguart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                 // jtaguart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> jtaguart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          jtaguart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;                       // jtaguart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> jtaguart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          jtaguart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;               // jtaguart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> jtaguart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [113:0] jtaguart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data;                        // jtaguart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> jtaguart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          jtaguart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;                       // jtaguart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> jtaguart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          jtaguart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;              // jtaguart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> jtaguart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          jtaguart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                    // jtaguart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> jtaguart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          jtaguart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;            // jtaguart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> jtaguart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [113:0] jtaguart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                     // jtaguart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> jtaguart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          jtaguart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                    // jtaguart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> jtaguart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          jtaguart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                  // jtaguart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> jtaguart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] jtaguart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                   // jtaguart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> jtaguart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          jtaguart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                  // jtaguart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> jtaguart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          prio_arbiter_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                   // prio_arbiter_0_s1_translator:uav_waitrequest -> prio_arbiter_0_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] prio_arbiter_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                    // prio_arbiter_0_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> prio_arbiter_0_s1_translator:uav_burstcount
	wire   [31:0] prio_arbiter_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                     // prio_arbiter_0_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> prio_arbiter_0_s1_translator:uav_writedata
	wire   [31:0] prio_arbiter_0_s1_translator_avalon_universal_slave_0_agent_m0_address;                                       // prio_arbiter_0_s1_translator_avalon_universal_slave_0_agent:m0_address -> prio_arbiter_0_s1_translator:uav_address
	wire          prio_arbiter_0_s1_translator_avalon_universal_slave_0_agent_m0_write;                                         // prio_arbiter_0_s1_translator_avalon_universal_slave_0_agent:m0_write -> prio_arbiter_0_s1_translator:uav_write
	wire          prio_arbiter_0_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                          // prio_arbiter_0_s1_translator_avalon_universal_slave_0_agent:m0_lock -> prio_arbiter_0_s1_translator:uav_lock
	wire          prio_arbiter_0_s1_translator_avalon_universal_slave_0_agent_m0_read;                                          // prio_arbiter_0_s1_translator_avalon_universal_slave_0_agent:m0_read -> prio_arbiter_0_s1_translator:uav_read
	wire   [31:0] prio_arbiter_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                      // prio_arbiter_0_s1_translator:uav_readdata -> prio_arbiter_0_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          prio_arbiter_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                 // prio_arbiter_0_s1_translator:uav_readdatavalid -> prio_arbiter_0_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          prio_arbiter_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                   // prio_arbiter_0_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> prio_arbiter_0_s1_translator:uav_debugaccess
	wire    [3:0] prio_arbiter_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                    // prio_arbiter_0_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> prio_arbiter_0_s1_translator:uav_byteenable
	wire          prio_arbiter_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                            // prio_arbiter_0_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> prio_arbiter_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          prio_arbiter_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                  // prio_arbiter_0_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> prio_arbiter_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          prio_arbiter_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                          // prio_arbiter_0_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> prio_arbiter_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [113:0] prio_arbiter_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                   // prio_arbiter_0_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> prio_arbiter_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          prio_arbiter_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                  // prio_arbiter_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> prio_arbiter_0_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          prio_arbiter_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                         // prio_arbiter_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> prio_arbiter_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          prio_arbiter_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                               // prio_arbiter_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> prio_arbiter_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          prio_arbiter_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                       // prio_arbiter_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> prio_arbiter_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [113:0] prio_arbiter_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                // prio_arbiter_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> prio_arbiter_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          prio_arbiter_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                               // prio_arbiter_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> prio_arbiter_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          prio_arbiter_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                             // prio_arbiter_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> prio_arbiter_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] prio_arbiter_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                              // prio_arbiter_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> prio_arbiter_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          prio_arbiter_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                             // prio_arbiter_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> prio_arbiter_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          traffic_gen_0_avalon_master_0_translator_avalon_universal_master_0_waitrequest;                               // traffic_gen_0_avalon_master_0_translator_avalon_universal_master_0_agent:av_waitrequest -> traffic_gen_0_avalon_master_0_translator:uav_waitrequest
	wire    [5:0] traffic_gen_0_avalon_master_0_translator_avalon_universal_master_0_burstcount;                                // traffic_gen_0_avalon_master_0_translator:uav_burstcount -> traffic_gen_0_avalon_master_0_translator_avalon_universal_master_0_agent:av_burstcount
	wire   [31:0] traffic_gen_0_avalon_master_0_translator_avalon_universal_master_0_writedata;                                 // traffic_gen_0_avalon_master_0_translator:uav_writedata -> traffic_gen_0_avalon_master_0_translator_avalon_universal_master_0_agent:av_writedata
	wire   [27:0] traffic_gen_0_avalon_master_0_translator_avalon_universal_master_0_address;                                   // traffic_gen_0_avalon_master_0_translator:uav_address -> traffic_gen_0_avalon_master_0_translator_avalon_universal_master_0_agent:av_address
	wire          traffic_gen_0_avalon_master_0_translator_avalon_universal_master_0_lock;                                      // traffic_gen_0_avalon_master_0_translator:uav_lock -> traffic_gen_0_avalon_master_0_translator_avalon_universal_master_0_agent:av_lock
	wire          traffic_gen_0_avalon_master_0_translator_avalon_universal_master_0_write;                                     // traffic_gen_0_avalon_master_0_translator:uav_write -> traffic_gen_0_avalon_master_0_translator_avalon_universal_master_0_agent:av_write
	wire          traffic_gen_0_avalon_master_0_translator_avalon_universal_master_0_read;                                      // traffic_gen_0_avalon_master_0_translator:uav_read -> traffic_gen_0_avalon_master_0_translator_avalon_universal_master_0_agent:av_read
	wire   [31:0] traffic_gen_0_avalon_master_0_translator_avalon_universal_master_0_readdata;                                  // traffic_gen_0_avalon_master_0_translator_avalon_universal_master_0_agent:av_readdata -> traffic_gen_0_avalon_master_0_translator:uav_readdata
	wire          traffic_gen_0_avalon_master_0_translator_avalon_universal_master_0_debugaccess;                               // traffic_gen_0_avalon_master_0_translator:uav_debugaccess -> traffic_gen_0_avalon_master_0_translator_avalon_universal_master_0_agent:av_debugaccess
	wire    [3:0] traffic_gen_0_avalon_master_0_translator_avalon_universal_master_0_byteenable;                                // traffic_gen_0_avalon_master_0_translator:uav_byteenable -> traffic_gen_0_avalon_master_0_translator_avalon_universal_master_0_agent:av_byteenable
	wire          traffic_gen_0_avalon_master_0_translator_avalon_universal_master_0_readdatavalid;                             // traffic_gen_0_avalon_master_0_translator_avalon_universal_master_0_agent:av_readdatavalid -> traffic_gen_0_avalon_master_0_translator:uav_readdatavalid
	wire          prio_arbiter_0_s2_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                   // prio_arbiter_0_s2_translator:uav_waitrequest -> prio_arbiter_0_s2_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] prio_arbiter_0_s2_translator_avalon_universal_slave_0_agent_m0_burstcount;                                    // prio_arbiter_0_s2_translator_avalon_universal_slave_0_agent:m0_burstcount -> prio_arbiter_0_s2_translator:uav_burstcount
	wire   [31:0] prio_arbiter_0_s2_translator_avalon_universal_slave_0_agent_m0_writedata;                                     // prio_arbiter_0_s2_translator_avalon_universal_slave_0_agent:m0_writedata -> prio_arbiter_0_s2_translator:uav_writedata
	wire   [27:0] prio_arbiter_0_s2_translator_avalon_universal_slave_0_agent_m0_address;                                       // prio_arbiter_0_s2_translator_avalon_universal_slave_0_agent:m0_address -> prio_arbiter_0_s2_translator:uav_address
	wire          prio_arbiter_0_s2_translator_avalon_universal_slave_0_agent_m0_write;                                         // prio_arbiter_0_s2_translator_avalon_universal_slave_0_agent:m0_write -> prio_arbiter_0_s2_translator:uav_write
	wire          prio_arbiter_0_s2_translator_avalon_universal_slave_0_agent_m0_lock;                                          // prio_arbiter_0_s2_translator_avalon_universal_slave_0_agent:m0_lock -> prio_arbiter_0_s2_translator:uav_lock
	wire          prio_arbiter_0_s2_translator_avalon_universal_slave_0_agent_m0_read;                                          // prio_arbiter_0_s2_translator_avalon_universal_slave_0_agent:m0_read -> prio_arbiter_0_s2_translator:uav_read
	wire   [31:0] prio_arbiter_0_s2_translator_avalon_universal_slave_0_agent_m0_readdata;                                      // prio_arbiter_0_s2_translator:uav_readdata -> prio_arbiter_0_s2_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          prio_arbiter_0_s2_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                 // prio_arbiter_0_s2_translator:uav_readdatavalid -> prio_arbiter_0_s2_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          prio_arbiter_0_s2_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                   // prio_arbiter_0_s2_translator_avalon_universal_slave_0_agent:m0_debugaccess -> prio_arbiter_0_s2_translator:uav_debugaccess
	wire    [3:0] prio_arbiter_0_s2_translator_avalon_universal_slave_0_agent_m0_byteenable;                                    // prio_arbiter_0_s2_translator_avalon_universal_slave_0_agent:m0_byteenable -> prio_arbiter_0_s2_translator:uav_byteenable
	wire          prio_arbiter_0_s2_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                            // prio_arbiter_0_s2_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> prio_arbiter_0_s2_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          prio_arbiter_0_s2_translator_avalon_universal_slave_0_agent_rf_source_valid;                                  // prio_arbiter_0_s2_translator_avalon_universal_slave_0_agent:rf_source_valid -> prio_arbiter_0_s2_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          prio_arbiter_0_s2_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                          // prio_arbiter_0_s2_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> prio_arbiter_0_s2_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [103:0] prio_arbiter_0_s2_translator_avalon_universal_slave_0_agent_rf_source_data;                                   // prio_arbiter_0_s2_translator_avalon_universal_slave_0_agent:rf_source_data -> prio_arbiter_0_s2_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          prio_arbiter_0_s2_translator_avalon_universal_slave_0_agent_rf_source_ready;                                  // prio_arbiter_0_s2_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> prio_arbiter_0_s2_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          prio_arbiter_0_s2_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                         // prio_arbiter_0_s2_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> prio_arbiter_0_s2_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          prio_arbiter_0_s2_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                               // prio_arbiter_0_s2_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> prio_arbiter_0_s2_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          prio_arbiter_0_s2_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                       // prio_arbiter_0_s2_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> prio_arbiter_0_s2_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [103:0] prio_arbiter_0_s2_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                // prio_arbiter_0_s2_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> prio_arbiter_0_s2_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          prio_arbiter_0_s2_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                               // prio_arbiter_0_s2_translator_avalon_universal_slave_0_agent:rf_sink_ready -> prio_arbiter_0_s2_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          prio_arbiter_0_s2_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                             // prio_arbiter_0_s2_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> prio_arbiter_0_s2_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] prio_arbiter_0_s2_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                              // prio_arbiter_0_s2_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> prio_arbiter_0_s2_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          prio_arbiter_0_s2_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                             // prio_arbiter_0_s2_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> prio_arbiter_0_s2_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          traffic_gen_1_avalon_master_0_translator_avalon_universal_master_0_waitrequest;                               // traffic_gen_1_avalon_master_0_translator_avalon_universal_master_0_agent:av_waitrequest -> traffic_gen_1_avalon_master_0_translator:uav_waitrequest
	wire    [5:0] traffic_gen_1_avalon_master_0_translator_avalon_universal_master_0_burstcount;                                // traffic_gen_1_avalon_master_0_translator:uav_burstcount -> traffic_gen_1_avalon_master_0_translator_avalon_universal_master_0_agent:av_burstcount
	wire   [31:0] traffic_gen_1_avalon_master_0_translator_avalon_universal_master_0_writedata;                                 // traffic_gen_1_avalon_master_0_translator:uav_writedata -> traffic_gen_1_avalon_master_0_translator_avalon_universal_master_0_agent:av_writedata
	wire   [27:0] traffic_gen_1_avalon_master_0_translator_avalon_universal_master_0_address;                                   // traffic_gen_1_avalon_master_0_translator:uav_address -> traffic_gen_1_avalon_master_0_translator_avalon_universal_master_0_agent:av_address
	wire          traffic_gen_1_avalon_master_0_translator_avalon_universal_master_0_lock;                                      // traffic_gen_1_avalon_master_0_translator:uav_lock -> traffic_gen_1_avalon_master_0_translator_avalon_universal_master_0_agent:av_lock
	wire          traffic_gen_1_avalon_master_0_translator_avalon_universal_master_0_write;                                     // traffic_gen_1_avalon_master_0_translator:uav_write -> traffic_gen_1_avalon_master_0_translator_avalon_universal_master_0_agent:av_write
	wire          traffic_gen_1_avalon_master_0_translator_avalon_universal_master_0_read;                                      // traffic_gen_1_avalon_master_0_translator:uav_read -> traffic_gen_1_avalon_master_0_translator_avalon_universal_master_0_agent:av_read
	wire   [31:0] traffic_gen_1_avalon_master_0_translator_avalon_universal_master_0_readdata;                                  // traffic_gen_1_avalon_master_0_translator_avalon_universal_master_0_agent:av_readdata -> traffic_gen_1_avalon_master_0_translator:uav_readdata
	wire          traffic_gen_1_avalon_master_0_translator_avalon_universal_master_0_debugaccess;                               // traffic_gen_1_avalon_master_0_translator:uav_debugaccess -> traffic_gen_1_avalon_master_0_translator_avalon_universal_master_0_agent:av_debugaccess
	wire    [3:0] traffic_gen_1_avalon_master_0_translator_avalon_universal_master_0_byteenable;                                // traffic_gen_1_avalon_master_0_translator:uav_byteenable -> traffic_gen_1_avalon_master_0_translator_avalon_universal_master_0_agent:av_byteenable
	wire          traffic_gen_1_avalon_master_0_translator_avalon_universal_master_0_readdatavalid;                             // traffic_gen_1_avalon_master_0_translator_avalon_universal_master_0_agent:av_readdatavalid -> traffic_gen_1_avalon_master_0_translator:uav_readdatavalid
	wire          prio_arbiter_0_s3_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                   // prio_arbiter_0_s3_translator:uav_waitrequest -> prio_arbiter_0_s3_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] prio_arbiter_0_s3_translator_avalon_universal_slave_0_agent_m0_burstcount;                                    // prio_arbiter_0_s3_translator_avalon_universal_slave_0_agent:m0_burstcount -> prio_arbiter_0_s3_translator:uav_burstcount
	wire   [31:0] prio_arbiter_0_s3_translator_avalon_universal_slave_0_agent_m0_writedata;                                     // prio_arbiter_0_s3_translator_avalon_universal_slave_0_agent:m0_writedata -> prio_arbiter_0_s3_translator:uav_writedata
	wire   [27:0] prio_arbiter_0_s3_translator_avalon_universal_slave_0_agent_m0_address;                                       // prio_arbiter_0_s3_translator_avalon_universal_slave_0_agent:m0_address -> prio_arbiter_0_s3_translator:uav_address
	wire          prio_arbiter_0_s3_translator_avalon_universal_slave_0_agent_m0_write;                                         // prio_arbiter_0_s3_translator_avalon_universal_slave_0_agent:m0_write -> prio_arbiter_0_s3_translator:uav_write
	wire          prio_arbiter_0_s3_translator_avalon_universal_slave_0_agent_m0_lock;                                          // prio_arbiter_0_s3_translator_avalon_universal_slave_0_agent:m0_lock -> prio_arbiter_0_s3_translator:uav_lock
	wire          prio_arbiter_0_s3_translator_avalon_universal_slave_0_agent_m0_read;                                          // prio_arbiter_0_s3_translator_avalon_universal_slave_0_agent:m0_read -> prio_arbiter_0_s3_translator:uav_read
	wire   [31:0] prio_arbiter_0_s3_translator_avalon_universal_slave_0_agent_m0_readdata;                                      // prio_arbiter_0_s3_translator:uav_readdata -> prio_arbiter_0_s3_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          prio_arbiter_0_s3_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                 // prio_arbiter_0_s3_translator:uav_readdatavalid -> prio_arbiter_0_s3_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          prio_arbiter_0_s3_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                   // prio_arbiter_0_s3_translator_avalon_universal_slave_0_agent:m0_debugaccess -> prio_arbiter_0_s3_translator:uav_debugaccess
	wire    [3:0] prio_arbiter_0_s3_translator_avalon_universal_slave_0_agent_m0_byteenable;                                    // prio_arbiter_0_s3_translator_avalon_universal_slave_0_agent:m0_byteenable -> prio_arbiter_0_s3_translator:uav_byteenable
	wire          prio_arbiter_0_s3_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                            // prio_arbiter_0_s3_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> prio_arbiter_0_s3_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          prio_arbiter_0_s3_translator_avalon_universal_slave_0_agent_rf_source_valid;                                  // prio_arbiter_0_s3_translator_avalon_universal_slave_0_agent:rf_source_valid -> prio_arbiter_0_s3_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          prio_arbiter_0_s3_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                          // prio_arbiter_0_s3_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> prio_arbiter_0_s3_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [103:0] prio_arbiter_0_s3_translator_avalon_universal_slave_0_agent_rf_source_data;                                   // prio_arbiter_0_s3_translator_avalon_universal_slave_0_agent:rf_source_data -> prio_arbiter_0_s3_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          prio_arbiter_0_s3_translator_avalon_universal_slave_0_agent_rf_source_ready;                                  // prio_arbiter_0_s3_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> prio_arbiter_0_s3_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          prio_arbiter_0_s3_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                         // prio_arbiter_0_s3_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> prio_arbiter_0_s3_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          prio_arbiter_0_s3_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                               // prio_arbiter_0_s3_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> prio_arbiter_0_s3_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          prio_arbiter_0_s3_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                       // prio_arbiter_0_s3_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> prio_arbiter_0_s3_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [103:0] prio_arbiter_0_s3_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                // prio_arbiter_0_s3_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> prio_arbiter_0_s3_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          prio_arbiter_0_s3_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                               // prio_arbiter_0_s3_translator_avalon_universal_slave_0_agent:rf_sink_ready -> prio_arbiter_0_s3_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          prio_arbiter_0_s3_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                             // prio_arbiter_0_s3_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> prio_arbiter_0_s3_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] prio_arbiter_0_s3_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                              // prio_arbiter_0_s3_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> prio_arbiter_0_s3_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          prio_arbiter_0_s3_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                             // prio_arbiter_0_s3_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> prio_arbiter_0_s3_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          com_nios_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket;                        // com_nios_instruction_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router:sink_endofpacket
	wire          com_nios_instruction_master_translator_avalon_universal_master_0_agent_cp_valid;                              // com_nios_instruction_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router:sink_valid
	wire          com_nios_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket;                      // com_nios_instruction_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router:sink_startofpacket
	wire  [112:0] com_nios_instruction_master_translator_avalon_universal_master_0_agent_cp_data;                               // com_nios_instruction_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router:sink_data
	wire          com_nios_instruction_master_translator_avalon_universal_master_0_agent_cp_ready;                              // addr_router:sink_ready -> com_nios_instruction_master_translator_avalon_universal_master_0_agent:cp_ready
	wire          com_nios_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket;                               // com_nios_data_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_001:sink_endofpacket
	wire          com_nios_data_master_translator_avalon_universal_master_0_agent_cp_valid;                                     // com_nios_data_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_001:sink_valid
	wire          com_nios_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket;                             // com_nios_data_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_001:sink_startofpacket
	wire  [112:0] com_nios_data_master_translator_avalon_universal_master_0_agent_cp_data;                                      // com_nios_data_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router_001:sink_data
	wire          com_nios_data_master_translator_avalon_universal_master_0_agent_cp_ready;                                     // addr_router_001:sink_ready -> com_nios_data_master_translator_avalon_universal_master_0_agent:cp_ready
	wire          carcontrol_nios_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket;                        // carControl_nios_data_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_002:sink_endofpacket
	wire          carcontrol_nios_data_master_translator_avalon_universal_master_0_agent_cp_valid;                              // carControl_nios_data_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_002:sink_valid
	wire          carcontrol_nios_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket;                      // carControl_nios_data_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_002:sink_startofpacket
	wire  [112:0] carcontrol_nios_data_master_translator_avalon_universal_master_0_agent_cp_data;                               // carControl_nios_data_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router_002:sink_data
	wire          carcontrol_nios_data_master_translator_avalon_universal_master_0_agent_cp_ready;                              // addr_router_002:sink_ready -> carControl_nios_data_master_translator_avalon_universal_master_0_agent:cp_ready
	wire          carcontrol_nios_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket;                 // carControl_nios_instruction_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_003:sink_endofpacket
	wire          carcontrol_nios_instruction_master_translator_avalon_universal_master_0_agent_cp_valid;                       // carControl_nios_instruction_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_003:sink_valid
	wire          carcontrol_nios_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket;               // carControl_nios_instruction_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_003:sink_startofpacket
	wire  [112:0] carcontrol_nios_instruction_master_translator_avalon_universal_master_0_agent_cp_data;                        // carControl_nios_instruction_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router_003:sink_data
	wire          carcontrol_nios_instruction_master_translator_avalon_universal_master_0_agent_cp_ready;                       // addr_router_003:sink_ready -> carControl_nios_instruction_master_translator_avalon_universal_master_0_agent:cp_ready
	wire          ethernet_subsystem_sgdma_rx_m_write_translator_avalon_universal_master_0_agent_cp_endofpacket;                // ethernet_subsystem_sgdma_rx_m_write_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_004:sink_endofpacket
	wire          ethernet_subsystem_sgdma_rx_m_write_translator_avalon_universal_master_0_agent_cp_valid;                      // ethernet_subsystem_sgdma_rx_m_write_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_004:sink_valid
	wire          ethernet_subsystem_sgdma_rx_m_write_translator_avalon_universal_master_0_agent_cp_startofpacket;              // ethernet_subsystem_sgdma_rx_m_write_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_004:sink_startofpacket
	wire  [112:0] ethernet_subsystem_sgdma_rx_m_write_translator_avalon_universal_master_0_agent_cp_data;                       // ethernet_subsystem_sgdma_rx_m_write_translator_avalon_universal_master_0_agent:cp_data -> addr_router_004:sink_data
	wire          ethernet_subsystem_sgdma_rx_m_write_translator_avalon_universal_master_0_agent_cp_ready;                      // addr_router_004:sink_ready -> ethernet_subsystem_sgdma_rx_m_write_translator_avalon_universal_master_0_agent:cp_ready
	wire          ethernet_subsystem_sgdma_tx_m_read_translator_avalon_universal_master_0_agent_cp_endofpacket;                 // ethernet_subsystem_sgdma_tx_m_read_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_005:sink_endofpacket
	wire          ethernet_subsystem_sgdma_tx_m_read_translator_avalon_universal_master_0_agent_cp_valid;                       // ethernet_subsystem_sgdma_tx_m_read_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_005:sink_valid
	wire          ethernet_subsystem_sgdma_tx_m_read_translator_avalon_universal_master_0_agent_cp_startofpacket;               // ethernet_subsystem_sgdma_tx_m_read_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_005:sink_startofpacket
	wire  [112:0] ethernet_subsystem_sgdma_tx_m_read_translator_avalon_universal_master_0_agent_cp_data;                        // ethernet_subsystem_sgdma_tx_m_read_translator_avalon_universal_master_0_agent:cp_data -> addr_router_005:sink_data
	wire          ethernet_subsystem_sgdma_tx_m_read_translator_avalon_universal_master_0_agent_cp_ready;                       // addr_router_005:sink_ready -> ethernet_subsystem_sgdma_tx_m_read_translator_avalon_universal_master_0_agent:cp_ready
	wire          com_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket;                          // com_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router:sink_endofpacket
	wire          com_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid;                                // com_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_valid -> id_router:sink_valid
	wire          com_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket;                        // com_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router:sink_startofpacket
	wire  [112:0] com_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data;                                 // com_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_data -> id_router:sink_data
	wire          com_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready;                                // id_router:sink_ready -> com_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_ready
	wire          com_memory_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                       // com_memory_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_001:sink_endofpacket
	wire          com_memory_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                             // com_memory_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_001:sink_valid
	wire          com_memory_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                     // com_memory_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_001:sink_startofpacket
	wire  [112:0] com_memory_s1_translator_avalon_universal_slave_0_agent_rp_data;                                              // com_memory_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_001:sink_data
	wire          com_memory_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                             // id_router_001:sink_ready -> com_memory_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          jtaguart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;                        // jtaguart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_002:sink_endofpacket
	wire          jtaguart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid;                              // jtaguart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_002:sink_valid
	wire          jtaguart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;                      // jtaguart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_002:sink_startofpacket
	wire  [112:0] jtaguart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data;                               // jtaguart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_002:sink_data
	wire          jtaguart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready;                              // id_router_002:sink_ready -> jtaguart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire          shared_memory_mutex_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                              // shared_memory_mutex_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_003:sink_endofpacket
	wire          shared_memory_mutex_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                    // shared_memory_mutex_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_003:sink_valid
	wire          shared_memory_mutex_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                            // shared_memory_mutex_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_003:sink_startofpacket
	wire  [112:0] shared_memory_mutex_s1_translator_avalon_universal_slave_0_agent_rp_data;                                     // shared_memory_mutex_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_003:sink_data
	wire          shared_memory_mutex_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                    // id_router_003:sink_ready -> shared_memory_mutex_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          com_timer_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                        // com_timer_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_004:sink_endofpacket
	wire          com_timer_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                              // com_timer_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_004:sink_valid
	wire          com_timer_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                      // com_timer_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_004:sink_startofpacket
	wire  [112:0] com_timer_s1_translator_avalon_universal_slave_0_agent_rp_data;                                               // com_timer_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_004:sink_data
	wire          com_timer_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                              // id_router_004:sink_ready -> com_timer_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          ethernet_subsystem_ethernet_bridge_s0_translator_avalon_universal_slave_0_agent_rp_endofpacket;               // ethernet_subsystem_ethernet_bridge_s0_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_005:sink_endofpacket
	wire          ethernet_subsystem_ethernet_bridge_s0_translator_avalon_universal_slave_0_agent_rp_valid;                     // ethernet_subsystem_ethernet_bridge_s0_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_005:sink_valid
	wire          ethernet_subsystem_ethernet_bridge_s0_translator_avalon_universal_slave_0_agent_rp_startofpacket;             // ethernet_subsystem_ethernet_bridge_s0_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_005:sink_startofpacket
	wire  [112:0] ethernet_subsystem_ethernet_bridge_s0_translator_avalon_universal_slave_0_agent_rp_data;                      // ethernet_subsystem_ethernet_bridge_s0_translator_avalon_universal_slave_0_agent:rp_data -> id_router_005:sink_data
	wire          ethernet_subsystem_ethernet_bridge_s0_translator_avalon_universal_slave_0_agent_rp_ready;                     // id_router_005:sink_ready -> ethernet_subsystem_ethernet_bridge_s0_translator_avalon_universal_slave_0_agent:rp_ready
	wire          ethernet_subsystem_descriptor_memory_s2_translator_avalon_universal_slave_0_agent_rp_endofpacket;             // ethernet_subsystem_descriptor_memory_s2_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_006:sink_endofpacket
	wire          ethernet_subsystem_descriptor_memory_s2_translator_avalon_universal_slave_0_agent_rp_valid;                   // ethernet_subsystem_descriptor_memory_s2_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_006:sink_valid
	wire          ethernet_subsystem_descriptor_memory_s2_translator_avalon_universal_slave_0_agent_rp_startofpacket;           // ethernet_subsystem_descriptor_memory_s2_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_006:sink_startofpacket
	wire  [112:0] ethernet_subsystem_descriptor_memory_s2_translator_avalon_universal_slave_0_agent_rp_data;                    // ethernet_subsystem_descriptor_memory_s2_translator_avalon_universal_slave_0_agent:rp_data -> id_router_006:sink_data
	wire          ethernet_subsystem_descriptor_memory_s2_translator_avalon_universal_slave_0_agent_rp_ready;                   // id_router_006:sink_ready -> ethernet_subsystem_descriptor_memory_s2_translator_avalon_universal_slave_0_agent:rp_ready
	wire          prio_arbiter_0_s0_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                   // prio_arbiter_0_s0_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_007:sink_endofpacket
	wire          prio_arbiter_0_s0_translator_avalon_universal_slave_0_agent_rp_valid;                                         // prio_arbiter_0_s0_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_007:sink_valid
	wire          prio_arbiter_0_s0_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                 // prio_arbiter_0_s0_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_007:sink_startofpacket
	wire  [112:0] prio_arbiter_0_s0_translator_avalon_universal_slave_0_agent_rp_data;                                          // prio_arbiter_0_s0_translator_avalon_universal_slave_0_agent:rp_data -> id_router_007:sink_data
	wire          prio_arbiter_0_s0_translator_avalon_universal_slave_0_agent_rp_ready;                                         // id_router_007:sink_ready -> prio_arbiter_0_s0_translator_avalon_universal_slave_0_agent:rp_ready
	wire          carcontrol_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket;                   // carControl_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_008:sink_endofpacket
	wire          carcontrol_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid;                         // carControl_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_008:sink_valid
	wire          carcontrol_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket;                 // carControl_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_008:sink_startofpacket
	wire  [112:0] carcontrol_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data;                          // carControl_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_data -> id_router_008:sink_data
	wire          carcontrol_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready;                         // id_router_008:sink_ready -> carControl_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_ready
	wire          onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                 // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_009:sink_endofpacket
	wire          onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                       // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_009:sink_valid
	wire          onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                               // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_009:sink_startofpacket
	wire  [112:0] onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rp_data;                                        // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_009:sink_data
	wire          onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                       // id_router_009:sink_ready -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          jtaguart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;                        // jtaguart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_010:sink_endofpacket
	wire          jtaguart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid;                              // jtaguart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_010:sink_valid
	wire          jtaguart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;                      // jtaguart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_010:sink_startofpacket
	wire  [112:0] jtaguart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data;                               // jtaguart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_010:sink_data
	wire          jtaguart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready;                              // id_router_010:sink_ready -> jtaguart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire          prio_arbiter_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                   // prio_arbiter_0_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_011:sink_endofpacket
	wire          prio_arbiter_0_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                         // prio_arbiter_0_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_011:sink_valid
	wire          prio_arbiter_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                 // prio_arbiter_0_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_011:sink_startofpacket
	wire  [112:0] prio_arbiter_0_s1_translator_avalon_universal_slave_0_agent_rp_data;                                          // prio_arbiter_0_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_011:sink_data
	wire          prio_arbiter_0_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                         // id_router_011:sink_ready -> prio_arbiter_0_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          traffic_gen_0_avalon_master_0_translator_avalon_universal_master_0_agent_cp_endofpacket;                      // traffic_gen_0_avalon_master_0_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_006:sink_endofpacket
	wire          traffic_gen_0_avalon_master_0_translator_avalon_universal_master_0_agent_cp_valid;                            // traffic_gen_0_avalon_master_0_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_006:sink_valid
	wire          traffic_gen_0_avalon_master_0_translator_avalon_universal_master_0_agent_cp_startofpacket;                    // traffic_gen_0_avalon_master_0_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_006:sink_startofpacket
	wire  [102:0] traffic_gen_0_avalon_master_0_translator_avalon_universal_master_0_agent_cp_data;                             // traffic_gen_0_avalon_master_0_translator_avalon_universal_master_0_agent:cp_data -> addr_router_006:sink_data
	wire          traffic_gen_0_avalon_master_0_translator_avalon_universal_master_0_agent_cp_ready;                            // addr_router_006:sink_ready -> traffic_gen_0_avalon_master_0_translator_avalon_universal_master_0_agent:cp_ready
	wire          prio_arbiter_0_s2_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                   // prio_arbiter_0_s2_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_012:sink_endofpacket
	wire          prio_arbiter_0_s2_translator_avalon_universal_slave_0_agent_rp_valid;                                         // prio_arbiter_0_s2_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_012:sink_valid
	wire          prio_arbiter_0_s2_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                 // prio_arbiter_0_s2_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_012:sink_startofpacket
	wire  [102:0] prio_arbiter_0_s2_translator_avalon_universal_slave_0_agent_rp_data;                                          // prio_arbiter_0_s2_translator_avalon_universal_slave_0_agent:rp_data -> id_router_012:sink_data
	wire          prio_arbiter_0_s2_translator_avalon_universal_slave_0_agent_rp_ready;                                         // id_router_012:sink_ready -> prio_arbiter_0_s2_translator_avalon_universal_slave_0_agent:rp_ready
	wire          traffic_gen_1_avalon_master_0_translator_avalon_universal_master_0_agent_cp_endofpacket;                      // traffic_gen_1_avalon_master_0_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_007:sink_endofpacket
	wire          traffic_gen_1_avalon_master_0_translator_avalon_universal_master_0_agent_cp_valid;                            // traffic_gen_1_avalon_master_0_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_007:sink_valid
	wire          traffic_gen_1_avalon_master_0_translator_avalon_universal_master_0_agent_cp_startofpacket;                    // traffic_gen_1_avalon_master_0_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_007:sink_startofpacket
	wire  [102:0] traffic_gen_1_avalon_master_0_translator_avalon_universal_master_0_agent_cp_data;                             // traffic_gen_1_avalon_master_0_translator_avalon_universal_master_0_agent:cp_data -> addr_router_007:sink_data
	wire          traffic_gen_1_avalon_master_0_translator_avalon_universal_master_0_agent_cp_ready;                            // addr_router_007:sink_ready -> traffic_gen_1_avalon_master_0_translator_avalon_universal_master_0_agent:cp_ready
	wire          prio_arbiter_0_s3_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                   // prio_arbiter_0_s3_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_013:sink_endofpacket
	wire          prio_arbiter_0_s3_translator_avalon_universal_slave_0_agent_rp_valid;                                         // prio_arbiter_0_s3_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_013:sink_valid
	wire          prio_arbiter_0_s3_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                 // prio_arbiter_0_s3_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_013:sink_startofpacket
	wire  [102:0] prio_arbiter_0_s3_translator_avalon_universal_slave_0_agent_rp_data;                                          // prio_arbiter_0_s3_translator_avalon_universal_slave_0_agent:rp_data -> id_router_013:sink_data
	wire          prio_arbiter_0_s3_translator_avalon_universal_slave_0_agent_rp_ready;                                         // id_router_013:sink_ready -> prio_arbiter_0_s3_translator_avalon_universal_slave_0_agent:rp_ready
	wire          addr_router_src_endofpacket;                                                                                  // addr_router:src_endofpacket -> limiter:cmd_sink_endofpacket
	wire          addr_router_src_valid;                                                                                        // addr_router:src_valid -> limiter:cmd_sink_valid
	wire          addr_router_src_startofpacket;                                                                                // addr_router:src_startofpacket -> limiter:cmd_sink_startofpacket
	wire  [112:0] addr_router_src_data;                                                                                         // addr_router:src_data -> limiter:cmd_sink_data
	wire   [11:0] addr_router_src_channel;                                                                                      // addr_router:src_channel -> limiter:cmd_sink_channel
	wire          addr_router_src_ready;                                                                                        // limiter:cmd_sink_ready -> addr_router:src_ready
	wire          limiter_rsp_src_endofpacket;                                                                                  // limiter:rsp_src_endofpacket -> com_nios_instruction_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire          limiter_rsp_src_valid;                                                                                        // limiter:rsp_src_valid -> com_nios_instruction_master_translator_avalon_universal_master_0_agent:rp_valid
	wire          limiter_rsp_src_startofpacket;                                                                                // limiter:rsp_src_startofpacket -> com_nios_instruction_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [112:0] limiter_rsp_src_data;                                                                                         // limiter:rsp_src_data -> com_nios_instruction_master_translator_avalon_universal_master_0_agent:rp_data
	wire   [11:0] limiter_rsp_src_channel;                                                                                      // limiter:rsp_src_channel -> com_nios_instruction_master_translator_avalon_universal_master_0_agent:rp_channel
	wire          limiter_rsp_src_ready;                                                                                        // com_nios_instruction_master_translator_avalon_universal_master_0_agent:rp_ready -> limiter:rsp_src_ready
	wire          addr_router_001_src_endofpacket;                                                                              // addr_router_001:src_endofpacket -> limiter_001:cmd_sink_endofpacket
	wire          addr_router_001_src_valid;                                                                                    // addr_router_001:src_valid -> limiter_001:cmd_sink_valid
	wire          addr_router_001_src_startofpacket;                                                                            // addr_router_001:src_startofpacket -> limiter_001:cmd_sink_startofpacket
	wire  [112:0] addr_router_001_src_data;                                                                                     // addr_router_001:src_data -> limiter_001:cmd_sink_data
	wire   [11:0] addr_router_001_src_channel;                                                                                  // addr_router_001:src_channel -> limiter_001:cmd_sink_channel
	wire          addr_router_001_src_ready;                                                                                    // limiter_001:cmd_sink_ready -> addr_router_001:src_ready
	wire          limiter_001_rsp_src_endofpacket;                                                                              // limiter_001:rsp_src_endofpacket -> com_nios_data_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire          limiter_001_rsp_src_valid;                                                                                    // limiter_001:rsp_src_valid -> com_nios_data_master_translator_avalon_universal_master_0_agent:rp_valid
	wire          limiter_001_rsp_src_startofpacket;                                                                            // limiter_001:rsp_src_startofpacket -> com_nios_data_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [112:0] limiter_001_rsp_src_data;                                                                                     // limiter_001:rsp_src_data -> com_nios_data_master_translator_avalon_universal_master_0_agent:rp_data
	wire   [11:0] limiter_001_rsp_src_channel;                                                                                  // limiter_001:rsp_src_channel -> com_nios_data_master_translator_avalon_universal_master_0_agent:rp_channel
	wire          limiter_001_rsp_src_ready;                                                                                    // com_nios_data_master_translator_avalon_universal_master_0_agent:rp_ready -> limiter_001:rsp_src_ready
	wire          addr_router_003_src_endofpacket;                                                                              // addr_router_003:src_endofpacket -> limiter_002:cmd_sink_endofpacket
	wire          addr_router_003_src_valid;                                                                                    // addr_router_003:src_valid -> limiter_002:cmd_sink_valid
	wire          addr_router_003_src_startofpacket;                                                                            // addr_router_003:src_startofpacket -> limiter_002:cmd_sink_startofpacket
	wire  [112:0] addr_router_003_src_data;                                                                                     // addr_router_003:src_data -> limiter_002:cmd_sink_data
	wire   [11:0] addr_router_003_src_channel;                                                                                  // addr_router_003:src_channel -> limiter_002:cmd_sink_channel
	wire          addr_router_003_src_ready;                                                                                    // limiter_002:cmd_sink_ready -> addr_router_003:src_ready
	wire          limiter_002_rsp_src_endofpacket;                                                                              // limiter_002:rsp_src_endofpacket -> carControl_nios_instruction_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire          limiter_002_rsp_src_valid;                                                                                    // limiter_002:rsp_src_valid -> carControl_nios_instruction_master_translator_avalon_universal_master_0_agent:rp_valid
	wire          limiter_002_rsp_src_startofpacket;                                                                            // limiter_002:rsp_src_startofpacket -> carControl_nios_instruction_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [112:0] limiter_002_rsp_src_data;                                                                                     // limiter_002:rsp_src_data -> carControl_nios_instruction_master_translator_avalon_universal_master_0_agent:rp_data
	wire   [11:0] limiter_002_rsp_src_channel;                                                                                  // limiter_002:rsp_src_channel -> carControl_nios_instruction_master_translator_avalon_universal_master_0_agent:rp_channel
	wire          limiter_002_rsp_src_ready;                                                                                    // carControl_nios_instruction_master_translator_avalon_universal_master_0_agent:rp_ready -> limiter_002:rsp_src_ready
	wire          burst_adapter_source0_endofpacket;                                                                            // burst_adapter:source0_endofpacket -> com_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          burst_adapter_source0_valid;                                                                                  // burst_adapter:source0_valid -> com_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_valid
	wire          burst_adapter_source0_startofpacket;                                                                          // burst_adapter:source0_startofpacket -> com_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [112:0] burst_adapter_source0_data;                                                                                   // burst_adapter:source0_data -> com_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_data
	wire          burst_adapter_source0_ready;                                                                                  // com_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter:source0_ready
	wire   [11:0] burst_adapter_source0_channel;                                                                                // burst_adapter:source0_channel -> com_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_channel
	wire          burst_adapter_001_source0_endofpacket;                                                                        // burst_adapter_001:source0_endofpacket -> com_memory_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          burst_adapter_001_source0_valid;                                                                              // burst_adapter_001:source0_valid -> com_memory_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          burst_adapter_001_source0_startofpacket;                                                                      // burst_adapter_001:source0_startofpacket -> com_memory_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [112:0] burst_adapter_001_source0_data;                                                                               // burst_adapter_001:source0_data -> com_memory_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire          burst_adapter_001_source0_ready;                                                                              // com_memory_s1_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter_001:source0_ready
	wire   [11:0] burst_adapter_001_source0_channel;                                                                            // burst_adapter_001:source0_channel -> com_memory_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          burst_adapter_002_source0_endofpacket;                                                                        // burst_adapter_002:source0_endofpacket -> jtaguart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          burst_adapter_002_source0_valid;                                                                              // burst_adapter_002:source0_valid -> jtaguart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire          burst_adapter_002_source0_startofpacket;                                                                      // burst_adapter_002:source0_startofpacket -> jtaguart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [112:0] burst_adapter_002_source0_data;                                                                               // burst_adapter_002:source0_data -> jtaguart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire          burst_adapter_002_source0_ready;                                                                              // jtaguart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter_002:source0_ready
	wire   [11:0] burst_adapter_002_source0_channel;                                                                            // burst_adapter_002:source0_channel -> jtaguart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire          burst_adapter_003_source0_endofpacket;                                                                        // burst_adapter_003:source0_endofpacket -> shared_memory_mutex_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          burst_adapter_003_source0_valid;                                                                              // burst_adapter_003:source0_valid -> shared_memory_mutex_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          burst_adapter_003_source0_startofpacket;                                                                      // burst_adapter_003:source0_startofpacket -> shared_memory_mutex_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [112:0] burst_adapter_003_source0_data;                                                                               // burst_adapter_003:source0_data -> shared_memory_mutex_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire          burst_adapter_003_source0_ready;                                                                              // shared_memory_mutex_s1_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter_003:source0_ready
	wire   [11:0] burst_adapter_003_source0_channel;                                                                            // burst_adapter_003:source0_channel -> shared_memory_mutex_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          burst_adapter_004_source0_endofpacket;                                                                        // burst_adapter_004:source0_endofpacket -> com_timer_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          burst_adapter_004_source0_valid;                                                                              // burst_adapter_004:source0_valid -> com_timer_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          burst_adapter_004_source0_startofpacket;                                                                      // burst_adapter_004:source0_startofpacket -> com_timer_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [112:0] burst_adapter_004_source0_data;                                                                               // burst_adapter_004:source0_data -> com_timer_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire          burst_adapter_004_source0_ready;                                                                              // com_timer_s1_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter_004:source0_ready
	wire   [11:0] burst_adapter_004_source0_channel;                                                                            // burst_adapter_004:source0_channel -> com_timer_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          burst_adapter_005_source0_endofpacket;                                                                        // burst_adapter_005:source0_endofpacket -> ethernet_subsystem_ethernet_bridge_s0_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          burst_adapter_005_source0_valid;                                                                              // burst_adapter_005:source0_valid -> ethernet_subsystem_ethernet_bridge_s0_translator_avalon_universal_slave_0_agent:cp_valid
	wire          burst_adapter_005_source0_startofpacket;                                                                      // burst_adapter_005:source0_startofpacket -> ethernet_subsystem_ethernet_bridge_s0_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [112:0] burst_adapter_005_source0_data;                                                                               // burst_adapter_005:source0_data -> ethernet_subsystem_ethernet_bridge_s0_translator_avalon_universal_slave_0_agent:cp_data
	wire          burst_adapter_005_source0_ready;                                                                              // ethernet_subsystem_ethernet_bridge_s0_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter_005:source0_ready
	wire   [11:0] burst_adapter_005_source0_channel;                                                                            // burst_adapter_005:source0_channel -> ethernet_subsystem_ethernet_bridge_s0_translator_avalon_universal_slave_0_agent:cp_channel
	wire          burst_adapter_006_source0_endofpacket;                                                                        // burst_adapter_006:source0_endofpacket -> ethernet_subsystem_descriptor_memory_s2_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          burst_adapter_006_source0_valid;                                                                              // burst_adapter_006:source0_valid -> ethernet_subsystem_descriptor_memory_s2_translator_avalon_universal_slave_0_agent:cp_valid
	wire          burst_adapter_006_source0_startofpacket;                                                                      // burst_adapter_006:source0_startofpacket -> ethernet_subsystem_descriptor_memory_s2_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [112:0] burst_adapter_006_source0_data;                                                                               // burst_adapter_006:source0_data -> ethernet_subsystem_descriptor_memory_s2_translator_avalon_universal_slave_0_agent:cp_data
	wire          burst_adapter_006_source0_ready;                                                                              // ethernet_subsystem_descriptor_memory_s2_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter_006:source0_ready
	wire   [11:0] burst_adapter_006_source0_channel;                                                                            // burst_adapter_006:source0_channel -> ethernet_subsystem_descriptor_memory_s2_translator_avalon_universal_slave_0_agent:cp_channel
	wire          burst_adapter_007_source0_endofpacket;                                                                        // burst_adapter_007:source0_endofpacket -> prio_arbiter_0_s0_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          burst_adapter_007_source0_valid;                                                                              // burst_adapter_007:source0_valid -> prio_arbiter_0_s0_translator_avalon_universal_slave_0_agent:cp_valid
	wire          burst_adapter_007_source0_startofpacket;                                                                      // burst_adapter_007:source0_startofpacket -> prio_arbiter_0_s0_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [112:0] burst_adapter_007_source0_data;                                                                               // burst_adapter_007:source0_data -> prio_arbiter_0_s0_translator_avalon_universal_slave_0_agent:cp_data
	wire          burst_adapter_007_source0_ready;                                                                              // prio_arbiter_0_s0_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter_007:source0_ready
	wire   [11:0] burst_adapter_007_source0_channel;                                                                            // burst_adapter_007:source0_channel -> prio_arbiter_0_s0_translator_avalon_universal_slave_0_agent:cp_channel
	wire          burst_adapter_008_source0_endofpacket;                                                                        // burst_adapter_008:source0_endofpacket -> prio_arbiter_0_s2_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          burst_adapter_008_source0_valid;                                                                              // burst_adapter_008:source0_valid -> prio_arbiter_0_s2_translator_avalon_universal_slave_0_agent:cp_valid
	wire          burst_adapter_008_source0_startofpacket;                                                                      // burst_adapter_008:source0_startofpacket -> prio_arbiter_0_s2_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [102:0] burst_adapter_008_source0_data;                                                                               // burst_adapter_008:source0_data -> prio_arbiter_0_s2_translator_avalon_universal_slave_0_agent:cp_data
	wire          burst_adapter_008_source0_ready;                                                                              // prio_arbiter_0_s2_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter_008:source0_ready
	wire          burst_adapter_008_source0_channel;                                                                            // burst_adapter_008:source0_channel -> prio_arbiter_0_s2_translator_avalon_universal_slave_0_agent:cp_channel
	wire          burst_adapter_009_source0_endofpacket;                                                                        // burst_adapter_009:source0_endofpacket -> prio_arbiter_0_s3_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          burst_adapter_009_source0_valid;                                                                              // burst_adapter_009:source0_valid -> prio_arbiter_0_s3_translator_avalon_universal_slave_0_agent:cp_valid
	wire          burst_adapter_009_source0_startofpacket;                                                                      // burst_adapter_009:source0_startofpacket -> prio_arbiter_0_s3_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [102:0] burst_adapter_009_source0_data;                                                                               // burst_adapter_009:source0_data -> prio_arbiter_0_s3_translator_avalon_universal_slave_0_agent:cp_data
	wire          burst_adapter_009_source0_ready;                                                                              // prio_arbiter_0_s3_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter_009:source0_ready
	wire          burst_adapter_009_source0_channel;                                                                            // burst_adapter_009:source0_channel -> prio_arbiter_0_s3_translator_avalon_universal_slave_0_agent:cp_channel
	wire          rst_controller_reset_out_reset;                                                                               // rst_controller:reset_out -> [addr_router:reset, addr_router_001:reset, addr_router_002:reset, addr_router_003:reset, addr_router_006:reset, addr_router_007:reset, burst_adapter:reset, burst_adapter_001:reset, burst_adapter_003:reset, burst_adapter_004:reset, burst_adapter_007:reset, burst_adapter_008:reset, burst_adapter_009:reset, carControl_nios:reset_n, carControl_nios_data_master_translator:reset, carControl_nios_data_master_translator_avalon_universal_master_0_agent:reset, carControl_nios_instruction_master_translator:reset, carControl_nios_instruction_master_translator_avalon_universal_master_0_agent:reset, carControl_nios_jtag_debug_module_translator:reset, carControl_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent:reset, carControl_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, cmd_xbar_demux:reset, cmd_xbar_demux_001:reset, cmd_xbar_demux_002:reset, cmd_xbar_demux_003:reset, cmd_xbar_demux_006:reset, cmd_xbar_demux_007:reset, cmd_xbar_mux:reset, cmd_xbar_mux_001:reset, cmd_xbar_mux_003:reset, cmd_xbar_mux_008:reset, cmd_xbar_mux_009:reset, com_memory:reset_n, com_memory_s1_translator:reset, com_memory_s1_translator_avalon_universal_slave_0_agent:reset, com_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, com_nios:reset_n, com_nios_data_master_translator:reset, com_nios_data_master_translator_avalon_universal_master_0_agent:reset, com_nios_instruction_master_translator:reset, com_nios_instruction_master_translator_avalon_universal_master_0_agent:reset, com_nios_jtag_debug_module_translator:reset, com_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent:reset, com_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, com_timer:reset_n, com_timer_s1_translator:reset, com_timer_s1_translator_avalon_universal_slave_0_agent:reset, com_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, id_router:reset, id_router_001:reset, id_router_003:reset, id_router_004:reset, id_router_007:reset, id_router_008:reset, id_router_009:reset, id_router_011:reset, id_router_012:reset, id_router_013:reset, irq_mapper:reset, irq_mapper_001:reset, limiter:reset, limiter_001:reset, limiter_002:reset, onchip_memory2_0:reset, onchip_memory2_0_s1_translator:reset, onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:reset, onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, prio_arbiter_0:csi_clockreset_RESET_n, prio_arbiter_0_m1_translator:reset, prio_arbiter_0_s0_translator:reset, prio_arbiter_0_s0_translator_avalon_universal_slave_0_agent:reset, prio_arbiter_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, prio_arbiter_0_s1_translator:reset, prio_arbiter_0_s1_translator_avalon_universal_slave_0_agent:reset, prio_arbiter_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, prio_arbiter_0_s2_translator:reset, prio_arbiter_0_s2_translator_avalon_universal_slave_0_agent:reset, prio_arbiter_0_s2_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, prio_arbiter_0_s3_translator:reset, prio_arbiter_0_s3_translator_avalon_universal_slave_0_agent:reset, prio_arbiter_0_s3_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, rsp_xbar_demux:reset, rsp_xbar_demux_001:reset, rsp_xbar_demux_003:reset, rsp_xbar_demux_004:reset, rsp_xbar_demux_007:reset, rsp_xbar_demux_008:reset, rsp_xbar_demux_009:reset, rsp_xbar_demux_011:reset, rsp_xbar_demux_012:reset, rsp_xbar_demux_013:reset, rsp_xbar_mux:reset, rsp_xbar_mux_001:reset, rsp_xbar_mux_002:reset, rsp_xbar_mux_003:reset, shared_memory:reset, shared_memory_mutex:reset_n, shared_memory_mutex_s1_translator:reset, shared_memory_mutex_s1_translator_avalon_universal_slave_0_agent:reset, shared_memory_mutex_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, shared_memory_s1_translator:reset, traffic_gen_0:iRESET, traffic_gen_0_avalon_master_0_translator:reset, traffic_gen_0_avalon_master_0_translator_avalon_universal_master_0_agent:reset, traffic_gen_1:iRESET, traffic_gen_1_avalon_master_0_translator:reset, traffic_gen_1_avalon_master_0_translator_avalon_universal_master_0_agent:reset]
	wire          com_nios_jtag_debug_module_reset_reset;                                                                       // com_nios:jtag_debug_module_resetrequest -> [rst_controller:reset_in1, rst_controller_001:reset_in1]
	wire          carcontrol_nios_jtag_debug_module_reset_reset;                                                                // carControl_nios:jtag_debug_module_resetrequest -> rst_controller:reset_in2
	wire          rst_controller_001_reset_out_reset;                                                                           // rst_controller_001:reset_out -> [burst_adapter_002:reset, id_router_002:reset, jtaguart_0:rst_n, jtaguart_0_avalon_jtag_slave_translator:reset, jtaguart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:reset, jtaguart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, rsp_xbar_demux_002:reset]
	wire          rst_controller_002_reset_out_reset;                                                                           // rst_controller_002:reset_out -> [addr_router_004:reset, addr_router_005:reset, burst_adapter_005:reset, burst_adapter_006:reset, cmd_xbar_demux_004:reset, cmd_xbar_demux_005:reset, ethernet_subsystem_descriptor_memory_s2_translator:reset, ethernet_subsystem_descriptor_memory_s2_translator_avalon_universal_slave_0_agent:reset, ethernet_subsystem_descriptor_memory_s2_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, ethernet_subsystem_ethernet_bridge_s0_translator:reset, ethernet_subsystem_ethernet_bridge_s0_translator_avalon_universal_slave_0_agent:reset, ethernet_subsystem_ethernet_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, ethernet_subsystem_sgdma_rx_m_write_translator:reset, ethernet_subsystem_sgdma_rx_m_write_translator_avalon_universal_master_0_agent:reset, ethernet_subsystem_sgdma_tx_m_read_translator:reset, ethernet_subsystem_sgdma_tx_m_read_translator_avalon_universal_master_0_agent:reset, id_router_005:reset, id_router_006:reset, id_router_010:reset, jtaguart_1:rst_n, jtaguart_1_avalon_jtag_slave_translator:reset, jtaguart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:reset, jtaguart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, rsp_xbar_demux_005:reset, rsp_xbar_demux_006:reset, rsp_xbar_demux_010:reset]
	wire          cmd_xbar_demux_src0_endofpacket;                                                                              // cmd_xbar_demux:src0_endofpacket -> cmd_xbar_mux:sink0_endofpacket
	wire          cmd_xbar_demux_src0_valid;                                                                                    // cmd_xbar_demux:src0_valid -> cmd_xbar_mux:sink0_valid
	wire          cmd_xbar_demux_src0_startofpacket;                                                                            // cmd_xbar_demux:src0_startofpacket -> cmd_xbar_mux:sink0_startofpacket
	wire  [112:0] cmd_xbar_demux_src0_data;                                                                                     // cmd_xbar_demux:src0_data -> cmd_xbar_mux:sink0_data
	wire   [11:0] cmd_xbar_demux_src0_channel;                                                                                  // cmd_xbar_demux:src0_channel -> cmd_xbar_mux:sink0_channel
	wire          cmd_xbar_demux_src0_ready;                                                                                    // cmd_xbar_mux:sink0_ready -> cmd_xbar_demux:src0_ready
	wire          cmd_xbar_demux_src1_endofpacket;                                                                              // cmd_xbar_demux:src1_endofpacket -> cmd_xbar_mux_001:sink0_endofpacket
	wire          cmd_xbar_demux_src1_valid;                                                                                    // cmd_xbar_demux:src1_valid -> cmd_xbar_mux_001:sink0_valid
	wire          cmd_xbar_demux_src1_startofpacket;                                                                            // cmd_xbar_demux:src1_startofpacket -> cmd_xbar_mux_001:sink0_startofpacket
	wire  [112:0] cmd_xbar_demux_src1_data;                                                                                     // cmd_xbar_demux:src1_data -> cmd_xbar_mux_001:sink0_data
	wire   [11:0] cmd_xbar_demux_src1_channel;                                                                                  // cmd_xbar_demux:src1_channel -> cmd_xbar_mux_001:sink0_channel
	wire          cmd_xbar_demux_src1_ready;                                                                                    // cmd_xbar_mux_001:sink0_ready -> cmd_xbar_demux:src1_ready
	wire          cmd_xbar_demux_001_src0_endofpacket;                                                                          // cmd_xbar_demux_001:src0_endofpacket -> cmd_xbar_mux:sink1_endofpacket
	wire          cmd_xbar_demux_001_src0_valid;                                                                                // cmd_xbar_demux_001:src0_valid -> cmd_xbar_mux:sink1_valid
	wire          cmd_xbar_demux_001_src0_startofpacket;                                                                        // cmd_xbar_demux_001:src0_startofpacket -> cmd_xbar_mux:sink1_startofpacket
	wire  [112:0] cmd_xbar_demux_001_src0_data;                                                                                 // cmd_xbar_demux_001:src0_data -> cmd_xbar_mux:sink1_data
	wire   [11:0] cmd_xbar_demux_001_src0_channel;                                                                              // cmd_xbar_demux_001:src0_channel -> cmd_xbar_mux:sink1_channel
	wire          cmd_xbar_demux_001_src0_ready;                                                                                // cmd_xbar_mux:sink1_ready -> cmd_xbar_demux_001:src0_ready
	wire          cmd_xbar_demux_001_src1_endofpacket;                                                                          // cmd_xbar_demux_001:src1_endofpacket -> cmd_xbar_mux_001:sink1_endofpacket
	wire          cmd_xbar_demux_001_src1_valid;                                                                                // cmd_xbar_demux_001:src1_valid -> cmd_xbar_mux_001:sink1_valid
	wire          cmd_xbar_demux_001_src1_startofpacket;                                                                        // cmd_xbar_demux_001:src1_startofpacket -> cmd_xbar_mux_001:sink1_startofpacket
	wire  [112:0] cmd_xbar_demux_001_src1_data;                                                                                 // cmd_xbar_demux_001:src1_data -> cmd_xbar_mux_001:sink1_data
	wire   [11:0] cmd_xbar_demux_001_src1_channel;                                                                              // cmd_xbar_demux_001:src1_channel -> cmd_xbar_mux_001:sink1_channel
	wire          cmd_xbar_demux_001_src1_ready;                                                                                // cmd_xbar_mux_001:sink1_ready -> cmd_xbar_demux_001:src1_ready
	wire          cmd_xbar_demux_001_src2_endofpacket;                                                                          // cmd_xbar_demux_001:src2_endofpacket -> burst_adapter_002:sink0_endofpacket
	wire          cmd_xbar_demux_001_src2_valid;                                                                                // cmd_xbar_demux_001:src2_valid -> burst_adapter_002:sink0_valid
	wire          cmd_xbar_demux_001_src2_startofpacket;                                                                        // cmd_xbar_demux_001:src2_startofpacket -> burst_adapter_002:sink0_startofpacket
	wire  [112:0] cmd_xbar_demux_001_src2_data;                                                                                 // cmd_xbar_demux_001:src2_data -> burst_adapter_002:sink0_data
	wire   [11:0] cmd_xbar_demux_001_src2_channel;                                                                              // cmd_xbar_demux_001:src2_channel -> burst_adapter_002:sink0_channel
	wire          cmd_xbar_demux_001_src3_endofpacket;                                                                          // cmd_xbar_demux_001:src3_endofpacket -> cmd_xbar_mux_003:sink0_endofpacket
	wire          cmd_xbar_demux_001_src3_valid;                                                                                // cmd_xbar_demux_001:src3_valid -> cmd_xbar_mux_003:sink0_valid
	wire          cmd_xbar_demux_001_src3_startofpacket;                                                                        // cmd_xbar_demux_001:src3_startofpacket -> cmd_xbar_mux_003:sink0_startofpacket
	wire  [112:0] cmd_xbar_demux_001_src3_data;                                                                                 // cmd_xbar_demux_001:src3_data -> cmd_xbar_mux_003:sink0_data
	wire   [11:0] cmd_xbar_demux_001_src3_channel;                                                                              // cmd_xbar_demux_001:src3_channel -> cmd_xbar_mux_003:sink0_channel
	wire          cmd_xbar_demux_001_src3_ready;                                                                                // cmd_xbar_mux_003:sink0_ready -> cmd_xbar_demux_001:src3_ready
	wire          cmd_xbar_demux_001_src4_endofpacket;                                                                          // cmd_xbar_demux_001:src4_endofpacket -> burst_adapter_004:sink0_endofpacket
	wire          cmd_xbar_demux_001_src4_valid;                                                                                // cmd_xbar_demux_001:src4_valid -> burst_adapter_004:sink0_valid
	wire          cmd_xbar_demux_001_src4_startofpacket;                                                                        // cmd_xbar_demux_001:src4_startofpacket -> burst_adapter_004:sink0_startofpacket
	wire  [112:0] cmd_xbar_demux_001_src4_data;                                                                                 // cmd_xbar_demux_001:src4_data -> burst_adapter_004:sink0_data
	wire   [11:0] cmd_xbar_demux_001_src4_channel;                                                                              // cmd_xbar_demux_001:src4_channel -> burst_adapter_004:sink0_channel
	wire          cmd_xbar_demux_001_src5_endofpacket;                                                                          // cmd_xbar_demux_001:src5_endofpacket -> burst_adapter_005:sink0_endofpacket
	wire          cmd_xbar_demux_001_src5_valid;                                                                                // cmd_xbar_demux_001:src5_valid -> burst_adapter_005:sink0_valid
	wire          cmd_xbar_demux_001_src5_startofpacket;                                                                        // cmd_xbar_demux_001:src5_startofpacket -> burst_adapter_005:sink0_startofpacket
	wire  [112:0] cmd_xbar_demux_001_src5_data;                                                                                 // cmd_xbar_demux_001:src5_data -> burst_adapter_005:sink0_data
	wire   [11:0] cmd_xbar_demux_001_src5_channel;                                                                              // cmd_xbar_demux_001:src5_channel -> burst_adapter_005:sink0_channel
	wire          cmd_xbar_demux_001_src6_endofpacket;                                                                          // cmd_xbar_demux_001:src6_endofpacket -> burst_adapter_006:sink0_endofpacket
	wire          cmd_xbar_demux_001_src6_valid;                                                                                // cmd_xbar_demux_001:src6_valid -> burst_adapter_006:sink0_valid
	wire          cmd_xbar_demux_001_src6_startofpacket;                                                                        // cmd_xbar_demux_001:src6_startofpacket -> burst_adapter_006:sink0_startofpacket
	wire  [112:0] cmd_xbar_demux_001_src6_data;                                                                                 // cmd_xbar_demux_001:src6_data -> burst_adapter_006:sink0_data
	wire   [11:0] cmd_xbar_demux_001_src6_channel;                                                                              // cmd_xbar_demux_001:src6_channel -> burst_adapter_006:sink0_channel
	wire          cmd_xbar_demux_001_src7_endofpacket;                                                                          // cmd_xbar_demux_001:src7_endofpacket -> burst_adapter_007:sink0_endofpacket
	wire          cmd_xbar_demux_001_src7_valid;                                                                                // cmd_xbar_demux_001:src7_valid -> burst_adapter_007:sink0_valid
	wire          cmd_xbar_demux_001_src7_startofpacket;                                                                        // cmd_xbar_demux_001:src7_startofpacket -> burst_adapter_007:sink0_startofpacket
	wire  [112:0] cmd_xbar_demux_001_src7_data;                                                                                 // cmd_xbar_demux_001:src7_data -> burst_adapter_007:sink0_data
	wire   [11:0] cmd_xbar_demux_001_src7_channel;                                                                              // cmd_xbar_demux_001:src7_channel -> burst_adapter_007:sink0_channel
	wire          cmd_xbar_demux_002_src0_endofpacket;                                                                          // cmd_xbar_demux_002:src0_endofpacket -> cmd_xbar_mux_003:sink1_endofpacket
	wire          cmd_xbar_demux_002_src0_valid;                                                                                // cmd_xbar_demux_002:src0_valid -> cmd_xbar_mux_003:sink1_valid
	wire          cmd_xbar_demux_002_src0_startofpacket;                                                                        // cmd_xbar_demux_002:src0_startofpacket -> cmd_xbar_mux_003:sink1_startofpacket
	wire  [112:0] cmd_xbar_demux_002_src0_data;                                                                                 // cmd_xbar_demux_002:src0_data -> cmd_xbar_mux_003:sink1_data
	wire   [11:0] cmd_xbar_demux_002_src0_channel;                                                                              // cmd_xbar_demux_002:src0_channel -> cmd_xbar_mux_003:sink1_channel
	wire          cmd_xbar_demux_002_src0_ready;                                                                                // cmd_xbar_mux_003:sink1_ready -> cmd_xbar_demux_002:src0_ready
	wire          cmd_xbar_demux_002_src1_endofpacket;                                                                          // cmd_xbar_demux_002:src1_endofpacket -> cmd_xbar_mux_008:sink0_endofpacket
	wire          cmd_xbar_demux_002_src1_valid;                                                                                // cmd_xbar_demux_002:src1_valid -> cmd_xbar_mux_008:sink0_valid
	wire          cmd_xbar_demux_002_src1_startofpacket;                                                                        // cmd_xbar_demux_002:src1_startofpacket -> cmd_xbar_mux_008:sink0_startofpacket
	wire  [112:0] cmd_xbar_demux_002_src1_data;                                                                                 // cmd_xbar_demux_002:src1_data -> cmd_xbar_mux_008:sink0_data
	wire   [11:0] cmd_xbar_demux_002_src1_channel;                                                                              // cmd_xbar_demux_002:src1_channel -> cmd_xbar_mux_008:sink0_channel
	wire          cmd_xbar_demux_002_src1_ready;                                                                                // cmd_xbar_mux_008:sink0_ready -> cmd_xbar_demux_002:src1_ready
	wire          cmd_xbar_demux_002_src2_endofpacket;                                                                          // cmd_xbar_demux_002:src2_endofpacket -> cmd_xbar_mux_009:sink0_endofpacket
	wire          cmd_xbar_demux_002_src2_valid;                                                                                // cmd_xbar_demux_002:src2_valid -> cmd_xbar_mux_009:sink0_valid
	wire          cmd_xbar_demux_002_src2_startofpacket;                                                                        // cmd_xbar_demux_002:src2_startofpacket -> cmd_xbar_mux_009:sink0_startofpacket
	wire  [112:0] cmd_xbar_demux_002_src2_data;                                                                                 // cmd_xbar_demux_002:src2_data -> cmd_xbar_mux_009:sink0_data
	wire   [11:0] cmd_xbar_demux_002_src2_channel;                                                                              // cmd_xbar_demux_002:src2_channel -> cmd_xbar_mux_009:sink0_channel
	wire          cmd_xbar_demux_002_src2_ready;                                                                                // cmd_xbar_mux_009:sink0_ready -> cmd_xbar_demux_002:src2_ready
	wire          cmd_xbar_demux_002_src3_endofpacket;                                                                          // cmd_xbar_demux_002:src3_endofpacket -> jtaguart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_002_src3_valid;                                                                                // cmd_xbar_demux_002:src3_valid -> jtaguart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_002_src3_startofpacket;                                                                        // cmd_xbar_demux_002:src3_startofpacket -> jtaguart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [112:0] cmd_xbar_demux_002_src3_data;                                                                                 // cmd_xbar_demux_002:src3_data -> jtaguart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire   [11:0] cmd_xbar_demux_002_src3_channel;                                                                              // cmd_xbar_demux_002:src3_channel -> jtaguart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_002_src4_endofpacket;                                                                          // cmd_xbar_demux_002:src4_endofpacket -> prio_arbiter_0_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_002_src4_valid;                                                                                // cmd_xbar_demux_002:src4_valid -> prio_arbiter_0_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_002_src4_startofpacket;                                                                        // cmd_xbar_demux_002:src4_startofpacket -> prio_arbiter_0_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [112:0] cmd_xbar_demux_002_src4_data;                                                                                 // cmd_xbar_demux_002:src4_data -> prio_arbiter_0_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [11:0] cmd_xbar_demux_002_src4_channel;                                                                              // cmd_xbar_demux_002:src4_channel -> prio_arbiter_0_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_003_src0_endofpacket;                                                                          // cmd_xbar_demux_003:src0_endofpacket -> cmd_xbar_mux_008:sink1_endofpacket
	wire          cmd_xbar_demux_003_src0_valid;                                                                                // cmd_xbar_demux_003:src0_valid -> cmd_xbar_mux_008:sink1_valid
	wire          cmd_xbar_demux_003_src0_startofpacket;                                                                        // cmd_xbar_demux_003:src0_startofpacket -> cmd_xbar_mux_008:sink1_startofpacket
	wire  [112:0] cmd_xbar_demux_003_src0_data;                                                                                 // cmd_xbar_demux_003:src0_data -> cmd_xbar_mux_008:sink1_data
	wire   [11:0] cmd_xbar_demux_003_src0_channel;                                                                              // cmd_xbar_demux_003:src0_channel -> cmd_xbar_mux_008:sink1_channel
	wire          cmd_xbar_demux_003_src0_ready;                                                                                // cmd_xbar_mux_008:sink1_ready -> cmd_xbar_demux_003:src0_ready
	wire          cmd_xbar_demux_003_src1_endofpacket;                                                                          // cmd_xbar_demux_003:src1_endofpacket -> cmd_xbar_mux_009:sink1_endofpacket
	wire          cmd_xbar_demux_003_src1_valid;                                                                                // cmd_xbar_demux_003:src1_valid -> cmd_xbar_mux_009:sink1_valid
	wire          cmd_xbar_demux_003_src1_startofpacket;                                                                        // cmd_xbar_demux_003:src1_startofpacket -> cmd_xbar_mux_009:sink1_startofpacket
	wire  [112:0] cmd_xbar_demux_003_src1_data;                                                                                 // cmd_xbar_demux_003:src1_data -> cmd_xbar_mux_009:sink1_data
	wire   [11:0] cmd_xbar_demux_003_src1_channel;                                                                              // cmd_xbar_demux_003:src1_channel -> cmd_xbar_mux_009:sink1_channel
	wire          cmd_xbar_demux_003_src1_ready;                                                                                // cmd_xbar_mux_009:sink1_ready -> cmd_xbar_demux_003:src1_ready
	wire          cmd_xbar_demux_004_src0_endofpacket;                                                                          // cmd_xbar_demux_004:src0_endofpacket -> cmd_xbar_mux_001:sink2_endofpacket
	wire          cmd_xbar_demux_004_src0_valid;                                                                                // cmd_xbar_demux_004:src0_valid -> cmd_xbar_mux_001:sink2_valid
	wire          cmd_xbar_demux_004_src0_startofpacket;                                                                        // cmd_xbar_demux_004:src0_startofpacket -> cmd_xbar_mux_001:sink2_startofpacket
	wire  [112:0] cmd_xbar_demux_004_src0_data;                                                                                 // cmd_xbar_demux_004:src0_data -> cmd_xbar_mux_001:sink2_data
	wire   [11:0] cmd_xbar_demux_004_src0_channel;                                                                              // cmd_xbar_demux_004:src0_channel -> cmd_xbar_mux_001:sink2_channel
	wire          cmd_xbar_demux_004_src0_ready;                                                                                // cmd_xbar_mux_001:sink2_ready -> cmd_xbar_demux_004:src0_ready
	wire          cmd_xbar_demux_005_src0_endofpacket;                                                                          // cmd_xbar_demux_005:src0_endofpacket -> cmd_xbar_mux_001:sink3_endofpacket
	wire          cmd_xbar_demux_005_src0_valid;                                                                                // cmd_xbar_demux_005:src0_valid -> cmd_xbar_mux_001:sink3_valid
	wire          cmd_xbar_demux_005_src0_startofpacket;                                                                        // cmd_xbar_demux_005:src0_startofpacket -> cmd_xbar_mux_001:sink3_startofpacket
	wire  [112:0] cmd_xbar_demux_005_src0_data;                                                                                 // cmd_xbar_demux_005:src0_data -> cmd_xbar_mux_001:sink3_data
	wire   [11:0] cmd_xbar_demux_005_src0_channel;                                                                              // cmd_xbar_demux_005:src0_channel -> cmd_xbar_mux_001:sink3_channel
	wire          cmd_xbar_demux_005_src0_ready;                                                                                // cmd_xbar_mux_001:sink3_ready -> cmd_xbar_demux_005:src0_ready
	wire          rsp_xbar_demux_src0_endofpacket;                                                                              // rsp_xbar_demux:src0_endofpacket -> rsp_xbar_mux:sink0_endofpacket
	wire          rsp_xbar_demux_src0_valid;                                                                                    // rsp_xbar_demux:src0_valid -> rsp_xbar_mux:sink0_valid
	wire          rsp_xbar_demux_src0_startofpacket;                                                                            // rsp_xbar_demux:src0_startofpacket -> rsp_xbar_mux:sink0_startofpacket
	wire  [112:0] rsp_xbar_demux_src0_data;                                                                                     // rsp_xbar_demux:src0_data -> rsp_xbar_mux:sink0_data
	wire   [11:0] rsp_xbar_demux_src0_channel;                                                                                  // rsp_xbar_demux:src0_channel -> rsp_xbar_mux:sink0_channel
	wire          rsp_xbar_demux_src0_ready;                                                                                    // rsp_xbar_mux:sink0_ready -> rsp_xbar_demux:src0_ready
	wire          rsp_xbar_demux_src1_endofpacket;                                                                              // rsp_xbar_demux:src1_endofpacket -> rsp_xbar_mux_001:sink0_endofpacket
	wire          rsp_xbar_demux_src1_valid;                                                                                    // rsp_xbar_demux:src1_valid -> rsp_xbar_mux_001:sink0_valid
	wire          rsp_xbar_demux_src1_startofpacket;                                                                            // rsp_xbar_demux:src1_startofpacket -> rsp_xbar_mux_001:sink0_startofpacket
	wire  [112:0] rsp_xbar_demux_src1_data;                                                                                     // rsp_xbar_demux:src1_data -> rsp_xbar_mux_001:sink0_data
	wire   [11:0] rsp_xbar_demux_src1_channel;                                                                                  // rsp_xbar_demux:src1_channel -> rsp_xbar_mux_001:sink0_channel
	wire          rsp_xbar_demux_src1_ready;                                                                                    // rsp_xbar_mux_001:sink0_ready -> rsp_xbar_demux:src1_ready
	wire          rsp_xbar_demux_001_src0_endofpacket;                                                                          // rsp_xbar_demux_001:src0_endofpacket -> rsp_xbar_mux:sink1_endofpacket
	wire          rsp_xbar_demux_001_src0_valid;                                                                                // rsp_xbar_demux_001:src0_valid -> rsp_xbar_mux:sink1_valid
	wire          rsp_xbar_demux_001_src0_startofpacket;                                                                        // rsp_xbar_demux_001:src0_startofpacket -> rsp_xbar_mux:sink1_startofpacket
	wire  [112:0] rsp_xbar_demux_001_src0_data;                                                                                 // rsp_xbar_demux_001:src0_data -> rsp_xbar_mux:sink1_data
	wire   [11:0] rsp_xbar_demux_001_src0_channel;                                                                              // rsp_xbar_demux_001:src0_channel -> rsp_xbar_mux:sink1_channel
	wire          rsp_xbar_demux_001_src0_ready;                                                                                // rsp_xbar_mux:sink1_ready -> rsp_xbar_demux_001:src0_ready
	wire          rsp_xbar_demux_001_src1_endofpacket;                                                                          // rsp_xbar_demux_001:src1_endofpacket -> rsp_xbar_mux_001:sink1_endofpacket
	wire          rsp_xbar_demux_001_src1_valid;                                                                                // rsp_xbar_demux_001:src1_valid -> rsp_xbar_mux_001:sink1_valid
	wire          rsp_xbar_demux_001_src1_startofpacket;                                                                        // rsp_xbar_demux_001:src1_startofpacket -> rsp_xbar_mux_001:sink1_startofpacket
	wire  [112:0] rsp_xbar_demux_001_src1_data;                                                                                 // rsp_xbar_demux_001:src1_data -> rsp_xbar_mux_001:sink1_data
	wire   [11:0] rsp_xbar_demux_001_src1_channel;                                                                              // rsp_xbar_demux_001:src1_channel -> rsp_xbar_mux_001:sink1_channel
	wire          rsp_xbar_demux_001_src1_ready;                                                                                // rsp_xbar_mux_001:sink1_ready -> rsp_xbar_demux_001:src1_ready
	wire          rsp_xbar_demux_001_src2_endofpacket;                                                                          // rsp_xbar_demux_001:src2_endofpacket -> ethernet_subsystem_sgdma_rx_m_write_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire          rsp_xbar_demux_001_src2_valid;                                                                                // rsp_xbar_demux_001:src2_valid -> ethernet_subsystem_sgdma_rx_m_write_translator_avalon_universal_master_0_agent:rp_valid
	wire          rsp_xbar_demux_001_src2_startofpacket;                                                                        // rsp_xbar_demux_001:src2_startofpacket -> ethernet_subsystem_sgdma_rx_m_write_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [112:0] rsp_xbar_demux_001_src2_data;                                                                                 // rsp_xbar_demux_001:src2_data -> ethernet_subsystem_sgdma_rx_m_write_translator_avalon_universal_master_0_agent:rp_data
	wire   [11:0] rsp_xbar_demux_001_src2_channel;                                                                              // rsp_xbar_demux_001:src2_channel -> ethernet_subsystem_sgdma_rx_m_write_translator_avalon_universal_master_0_agent:rp_channel
	wire          rsp_xbar_demux_001_src3_endofpacket;                                                                          // rsp_xbar_demux_001:src3_endofpacket -> ethernet_subsystem_sgdma_tx_m_read_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire          rsp_xbar_demux_001_src3_valid;                                                                                // rsp_xbar_demux_001:src3_valid -> ethernet_subsystem_sgdma_tx_m_read_translator_avalon_universal_master_0_agent:rp_valid
	wire          rsp_xbar_demux_001_src3_startofpacket;                                                                        // rsp_xbar_demux_001:src3_startofpacket -> ethernet_subsystem_sgdma_tx_m_read_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [112:0] rsp_xbar_demux_001_src3_data;                                                                                 // rsp_xbar_demux_001:src3_data -> ethernet_subsystem_sgdma_tx_m_read_translator_avalon_universal_master_0_agent:rp_data
	wire   [11:0] rsp_xbar_demux_001_src3_channel;                                                                              // rsp_xbar_demux_001:src3_channel -> ethernet_subsystem_sgdma_tx_m_read_translator_avalon_universal_master_0_agent:rp_channel
	wire          rsp_xbar_demux_002_src0_endofpacket;                                                                          // rsp_xbar_demux_002:src0_endofpacket -> rsp_xbar_mux_001:sink2_endofpacket
	wire          rsp_xbar_demux_002_src0_valid;                                                                                // rsp_xbar_demux_002:src0_valid -> rsp_xbar_mux_001:sink2_valid
	wire          rsp_xbar_demux_002_src0_startofpacket;                                                                        // rsp_xbar_demux_002:src0_startofpacket -> rsp_xbar_mux_001:sink2_startofpacket
	wire  [112:0] rsp_xbar_demux_002_src0_data;                                                                                 // rsp_xbar_demux_002:src0_data -> rsp_xbar_mux_001:sink2_data
	wire   [11:0] rsp_xbar_demux_002_src0_channel;                                                                              // rsp_xbar_demux_002:src0_channel -> rsp_xbar_mux_001:sink2_channel
	wire          rsp_xbar_demux_002_src0_ready;                                                                                // rsp_xbar_mux_001:sink2_ready -> rsp_xbar_demux_002:src0_ready
	wire          rsp_xbar_demux_003_src0_endofpacket;                                                                          // rsp_xbar_demux_003:src0_endofpacket -> rsp_xbar_mux_001:sink3_endofpacket
	wire          rsp_xbar_demux_003_src0_valid;                                                                                // rsp_xbar_demux_003:src0_valid -> rsp_xbar_mux_001:sink3_valid
	wire          rsp_xbar_demux_003_src0_startofpacket;                                                                        // rsp_xbar_demux_003:src0_startofpacket -> rsp_xbar_mux_001:sink3_startofpacket
	wire  [112:0] rsp_xbar_demux_003_src0_data;                                                                                 // rsp_xbar_demux_003:src0_data -> rsp_xbar_mux_001:sink3_data
	wire   [11:0] rsp_xbar_demux_003_src0_channel;                                                                              // rsp_xbar_demux_003:src0_channel -> rsp_xbar_mux_001:sink3_channel
	wire          rsp_xbar_demux_003_src0_ready;                                                                                // rsp_xbar_mux_001:sink3_ready -> rsp_xbar_demux_003:src0_ready
	wire          rsp_xbar_demux_003_src1_endofpacket;                                                                          // rsp_xbar_demux_003:src1_endofpacket -> rsp_xbar_mux_002:sink0_endofpacket
	wire          rsp_xbar_demux_003_src1_valid;                                                                                // rsp_xbar_demux_003:src1_valid -> rsp_xbar_mux_002:sink0_valid
	wire          rsp_xbar_demux_003_src1_startofpacket;                                                                        // rsp_xbar_demux_003:src1_startofpacket -> rsp_xbar_mux_002:sink0_startofpacket
	wire  [112:0] rsp_xbar_demux_003_src1_data;                                                                                 // rsp_xbar_demux_003:src1_data -> rsp_xbar_mux_002:sink0_data
	wire   [11:0] rsp_xbar_demux_003_src1_channel;                                                                              // rsp_xbar_demux_003:src1_channel -> rsp_xbar_mux_002:sink0_channel
	wire          rsp_xbar_demux_003_src1_ready;                                                                                // rsp_xbar_mux_002:sink0_ready -> rsp_xbar_demux_003:src1_ready
	wire          rsp_xbar_demux_004_src0_endofpacket;                                                                          // rsp_xbar_demux_004:src0_endofpacket -> rsp_xbar_mux_001:sink4_endofpacket
	wire          rsp_xbar_demux_004_src0_valid;                                                                                // rsp_xbar_demux_004:src0_valid -> rsp_xbar_mux_001:sink4_valid
	wire          rsp_xbar_demux_004_src0_startofpacket;                                                                        // rsp_xbar_demux_004:src0_startofpacket -> rsp_xbar_mux_001:sink4_startofpacket
	wire  [112:0] rsp_xbar_demux_004_src0_data;                                                                                 // rsp_xbar_demux_004:src0_data -> rsp_xbar_mux_001:sink4_data
	wire   [11:0] rsp_xbar_demux_004_src0_channel;                                                                              // rsp_xbar_demux_004:src0_channel -> rsp_xbar_mux_001:sink4_channel
	wire          rsp_xbar_demux_004_src0_ready;                                                                                // rsp_xbar_mux_001:sink4_ready -> rsp_xbar_demux_004:src0_ready
	wire          rsp_xbar_demux_005_src0_endofpacket;                                                                          // rsp_xbar_demux_005:src0_endofpacket -> rsp_xbar_mux_001:sink5_endofpacket
	wire          rsp_xbar_demux_005_src0_valid;                                                                                // rsp_xbar_demux_005:src0_valid -> rsp_xbar_mux_001:sink5_valid
	wire          rsp_xbar_demux_005_src0_startofpacket;                                                                        // rsp_xbar_demux_005:src0_startofpacket -> rsp_xbar_mux_001:sink5_startofpacket
	wire  [112:0] rsp_xbar_demux_005_src0_data;                                                                                 // rsp_xbar_demux_005:src0_data -> rsp_xbar_mux_001:sink5_data
	wire   [11:0] rsp_xbar_demux_005_src0_channel;                                                                              // rsp_xbar_demux_005:src0_channel -> rsp_xbar_mux_001:sink5_channel
	wire          rsp_xbar_demux_005_src0_ready;                                                                                // rsp_xbar_mux_001:sink5_ready -> rsp_xbar_demux_005:src0_ready
	wire          rsp_xbar_demux_006_src0_endofpacket;                                                                          // rsp_xbar_demux_006:src0_endofpacket -> rsp_xbar_mux_001:sink6_endofpacket
	wire          rsp_xbar_demux_006_src0_valid;                                                                                // rsp_xbar_demux_006:src0_valid -> rsp_xbar_mux_001:sink6_valid
	wire          rsp_xbar_demux_006_src0_startofpacket;                                                                        // rsp_xbar_demux_006:src0_startofpacket -> rsp_xbar_mux_001:sink6_startofpacket
	wire  [112:0] rsp_xbar_demux_006_src0_data;                                                                                 // rsp_xbar_demux_006:src0_data -> rsp_xbar_mux_001:sink6_data
	wire   [11:0] rsp_xbar_demux_006_src0_channel;                                                                              // rsp_xbar_demux_006:src0_channel -> rsp_xbar_mux_001:sink6_channel
	wire          rsp_xbar_demux_006_src0_ready;                                                                                // rsp_xbar_mux_001:sink6_ready -> rsp_xbar_demux_006:src0_ready
	wire          rsp_xbar_demux_007_src0_endofpacket;                                                                          // rsp_xbar_demux_007:src0_endofpacket -> rsp_xbar_mux_001:sink7_endofpacket
	wire          rsp_xbar_demux_007_src0_valid;                                                                                // rsp_xbar_demux_007:src0_valid -> rsp_xbar_mux_001:sink7_valid
	wire          rsp_xbar_demux_007_src0_startofpacket;                                                                        // rsp_xbar_demux_007:src0_startofpacket -> rsp_xbar_mux_001:sink7_startofpacket
	wire  [112:0] rsp_xbar_demux_007_src0_data;                                                                                 // rsp_xbar_demux_007:src0_data -> rsp_xbar_mux_001:sink7_data
	wire   [11:0] rsp_xbar_demux_007_src0_channel;                                                                              // rsp_xbar_demux_007:src0_channel -> rsp_xbar_mux_001:sink7_channel
	wire          rsp_xbar_demux_007_src0_ready;                                                                                // rsp_xbar_mux_001:sink7_ready -> rsp_xbar_demux_007:src0_ready
	wire          rsp_xbar_demux_008_src0_endofpacket;                                                                          // rsp_xbar_demux_008:src0_endofpacket -> rsp_xbar_mux_002:sink1_endofpacket
	wire          rsp_xbar_demux_008_src0_valid;                                                                                // rsp_xbar_demux_008:src0_valid -> rsp_xbar_mux_002:sink1_valid
	wire          rsp_xbar_demux_008_src0_startofpacket;                                                                        // rsp_xbar_demux_008:src0_startofpacket -> rsp_xbar_mux_002:sink1_startofpacket
	wire  [112:0] rsp_xbar_demux_008_src0_data;                                                                                 // rsp_xbar_demux_008:src0_data -> rsp_xbar_mux_002:sink1_data
	wire   [11:0] rsp_xbar_demux_008_src0_channel;                                                                              // rsp_xbar_demux_008:src0_channel -> rsp_xbar_mux_002:sink1_channel
	wire          rsp_xbar_demux_008_src0_ready;                                                                                // rsp_xbar_mux_002:sink1_ready -> rsp_xbar_demux_008:src0_ready
	wire          rsp_xbar_demux_008_src1_endofpacket;                                                                          // rsp_xbar_demux_008:src1_endofpacket -> rsp_xbar_mux_003:sink0_endofpacket
	wire          rsp_xbar_demux_008_src1_valid;                                                                                // rsp_xbar_demux_008:src1_valid -> rsp_xbar_mux_003:sink0_valid
	wire          rsp_xbar_demux_008_src1_startofpacket;                                                                        // rsp_xbar_demux_008:src1_startofpacket -> rsp_xbar_mux_003:sink0_startofpacket
	wire  [112:0] rsp_xbar_demux_008_src1_data;                                                                                 // rsp_xbar_demux_008:src1_data -> rsp_xbar_mux_003:sink0_data
	wire   [11:0] rsp_xbar_demux_008_src1_channel;                                                                              // rsp_xbar_demux_008:src1_channel -> rsp_xbar_mux_003:sink0_channel
	wire          rsp_xbar_demux_008_src1_ready;                                                                                // rsp_xbar_mux_003:sink0_ready -> rsp_xbar_demux_008:src1_ready
	wire          rsp_xbar_demux_009_src0_endofpacket;                                                                          // rsp_xbar_demux_009:src0_endofpacket -> rsp_xbar_mux_002:sink2_endofpacket
	wire          rsp_xbar_demux_009_src0_valid;                                                                                // rsp_xbar_demux_009:src0_valid -> rsp_xbar_mux_002:sink2_valid
	wire          rsp_xbar_demux_009_src0_startofpacket;                                                                        // rsp_xbar_demux_009:src0_startofpacket -> rsp_xbar_mux_002:sink2_startofpacket
	wire  [112:0] rsp_xbar_demux_009_src0_data;                                                                                 // rsp_xbar_demux_009:src0_data -> rsp_xbar_mux_002:sink2_data
	wire   [11:0] rsp_xbar_demux_009_src0_channel;                                                                              // rsp_xbar_demux_009:src0_channel -> rsp_xbar_mux_002:sink2_channel
	wire          rsp_xbar_demux_009_src0_ready;                                                                                // rsp_xbar_mux_002:sink2_ready -> rsp_xbar_demux_009:src0_ready
	wire          rsp_xbar_demux_009_src1_endofpacket;                                                                          // rsp_xbar_demux_009:src1_endofpacket -> rsp_xbar_mux_003:sink1_endofpacket
	wire          rsp_xbar_demux_009_src1_valid;                                                                                // rsp_xbar_demux_009:src1_valid -> rsp_xbar_mux_003:sink1_valid
	wire          rsp_xbar_demux_009_src1_startofpacket;                                                                        // rsp_xbar_demux_009:src1_startofpacket -> rsp_xbar_mux_003:sink1_startofpacket
	wire  [112:0] rsp_xbar_demux_009_src1_data;                                                                                 // rsp_xbar_demux_009:src1_data -> rsp_xbar_mux_003:sink1_data
	wire   [11:0] rsp_xbar_demux_009_src1_channel;                                                                              // rsp_xbar_demux_009:src1_channel -> rsp_xbar_mux_003:sink1_channel
	wire          rsp_xbar_demux_009_src1_ready;                                                                                // rsp_xbar_mux_003:sink1_ready -> rsp_xbar_demux_009:src1_ready
	wire          rsp_xbar_demux_010_src0_endofpacket;                                                                          // rsp_xbar_demux_010:src0_endofpacket -> rsp_xbar_mux_002:sink3_endofpacket
	wire          rsp_xbar_demux_010_src0_valid;                                                                                // rsp_xbar_demux_010:src0_valid -> rsp_xbar_mux_002:sink3_valid
	wire          rsp_xbar_demux_010_src0_startofpacket;                                                                        // rsp_xbar_demux_010:src0_startofpacket -> rsp_xbar_mux_002:sink3_startofpacket
	wire  [112:0] rsp_xbar_demux_010_src0_data;                                                                                 // rsp_xbar_demux_010:src0_data -> rsp_xbar_mux_002:sink3_data
	wire   [11:0] rsp_xbar_demux_010_src0_channel;                                                                              // rsp_xbar_demux_010:src0_channel -> rsp_xbar_mux_002:sink3_channel
	wire          rsp_xbar_demux_010_src0_ready;                                                                                // rsp_xbar_mux_002:sink3_ready -> rsp_xbar_demux_010:src0_ready
	wire          rsp_xbar_demux_011_src0_endofpacket;                                                                          // rsp_xbar_demux_011:src0_endofpacket -> rsp_xbar_mux_002:sink4_endofpacket
	wire          rsp_xbar_demux_011_src0_valid;                                                                                // rsp_xbar_demux_011:src0_valid -> rsp_xbar_mux_002:sink4_valid
	wire          rsp_xbar_demux_011_src0_startofpacket;                                                                        // rsp_xbar_demux_011:src0_startofpacket -> rsp_xbar_mux_002:sink4_startofpacket
	wire  [112:0] rsp_xbar_demux_011_src0_data;                                                                                 // rsp_xbar_demux_011:src0_data -> rsp_xbar_mux_002:sink4_data
	wire   [11:0] rsp_xbar_demux_011_src0_channel;                                                                              // rsp_xbar_demux_011:src0_channel -> rsp_xbar_mux_002:sink4_channel
	wire          rsp_xbar_demux_011_src0_ready;                                                                                // rsp_xbar_mux_002:sink4_ready -> rsp_xbar_demux_011:src0_ready
	wire          limiter_cmd_src_endofpacket;                                                                                  // limiter:cmd_src_endofpacket -> cmd_xbar_demux:sink_endofpacket
	wire          limiter_cmd_src_startofpacket;                                                                                // limiter:cmd_src_startofpacket -> cmd_xbar_demux:sink_startofpacket
	wire  [112:0] limiter_cmd_src_data;                                                                                         // limiter:cmd_src_data -> cmd_xbar_demux:sink_data
	wire   [11:0] limiter_cmd_src_channel;                                                                                      // limiter:cmd_src_channel -> cmd_xbar_demux:sink_channel
	wire          limiter_cmd_src_ready;                                                                                        // cmd_xbar_demux:sink_ready -> limiter:cmd_src_ready
	wire          rsp_xbar_mux_src_endofpacket;                                                                                 // rsp_xbar_mux:src_endofpacket -> limiter:rsp_sink_endofpacket
	wire          rsp_xbar_mux_src_valid;                                                                                       // rsp_xbar_mux:src_valid -> limiter:rsp_sink_valid
	wire          rsp_xbar_mux_src_startofpacket;                                                                               // rsp_xbar_mux:src_startofpacket -> limiter:rsp_sink_startofpacket
	wire  [112:0] rsp_xbar_mux_src_data;                                                                                        // rsp_xbar_mux:src_data -> limiter:rsp_sink_data
	wire   [11:0] rsp_xbar_mux_src_channel;                                                                                     // rsp_xbar_mux:src_channel -> limiter:rsp_sink_channel
	wire          rsp_xbar_mux_src_ready;                                                                                       // limiter:rsp_sink_ready -> rsp_xbar_mux:src_ready
	wire          limiter_001_cmd_src_endofpacket;                                                                              // limiter_001:cmd_src_endofpacket -> cmd_xbar_demux_001:sink_endofpacket
	wire          limiter_001_cmd_src_startofpacket;                                                                            // limiter_001:cmd_src_startofpacket -> cmd_xbar_demux_001:sink_startofpacket
	wire  [112:0] limiter_001_cmd_src_data;                                                                                     // limiter_001:cmd_src_data -> cmd_xbar_demux_001:sink_data
	wire   [11:0] limiter_001_cmd_src_channel;                                                                                  // limiter_001:cmd_src_channel -> cmd_xbar_demux_001:sink_channel
	wire          limiter_001_cmd_src_ready;                                                                                    // cmd_xbar_demux_001:sink_ready -> limiter_001:cmd_src_ready
	wire          rsp_xbar_mux_001_src_endofpacket;                                                                             // rsp_xbar_mux_001:src_endofpacket -> limiter_001:rsp_sink_endofpacket
	wire          rsp_xbar_mux_001_src_valid;                                                                                   // rsp_xbar_mux_001:src_valid -> limiter_001:rsp_sink_valid
	wire          rsp_xbar_mux_001_src_startofpacket;                                                                           // rsp_xbar_mux_001:src_startofpacket -> limiter_001:rsp_sink_startofpacket
	wire  [112:0] rsp_xbar_mux_001_src_data;                                                                                    // rsp_xbar_mux_001:src_data -> limiter_001:rsp_sink_data
	wire   [11:0] rsp_xbar_mux_001_src_channel;                                                                                 // rsp_xbar_mux_001:src_channel -> limiter_001:rsp_sink_channel
	wire          rsp_xbar_mux_001_src_ready;                                                                                   // limiter_001:rsp_sink_ready -> rsp_xbar_mux_001:src_ready
	wire          addr_router_002_src_endofpacket;                                                                              // addr_router_002:src_endofpacket -> cmd_xbar_demux_002:sink_endofpacket
	wire          addr_router_002_src_valid;                                                                                    // addr_router_002:src_valid -> cmd_xbar_demux_002:sink_valid
	wire          addr_router_002_src_startofpacket;                                                                            // addr_router_002:src_startofpacket -> cmd_xbar_demux_002:sink_startofpacket
	wire  [112:0] addr_router_002_src_data;                                                                                     // addr_router_002:src_data -> cmd_xbar_demux_002:sink_data
	wire   [11:0] addr_router_002_src_channel;                                                                                  // addr_router_002:src_channel -> cmd_xbar_demux_002:sink_channel
	wire          addr_router_002_src_ready;                                                                                    // cmd_xbar_demux_002:sink_ready -> addr_router_002:src_ready
	wire          rsp_xbar_mux_002_src_endofpacket;                                                                             // rsp_xbar_mux_002:src_endofpacket -> carControl_nios_data_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire          rsp_xbar_mux_002_src_valid;                                                                                   // rsp_xbar_mux_002:src_valid -> carControl_nios_data_master_translator_avalon_universal_master_0_agent:rp_valid
	wire          rsp_xbar_mux_002_src_startofpacket;                                                                           // rsp_xbar_mux_002:src_startofpacket -> carControl_nios_data_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [112:0] rsp_xbar_mux_002_src_data;                                                                                    // rsp_xbar_mux_002:src_data -> carControl_nios_data_master_translator_avalon_universal_master_0_agent:rp_data
	wire   [11:0] rsp_xbar_mux_002_src_channel;                                                                                 // rsp_xbar_mux_002:src_channel -> carControl_nios_data_master_translator_avalon_universal_master_0_agent:rp_channel
	wire          rsp_xbar_mux_002_src_ready;                                                                                   // carControl_nios_data_master_translator_avalon_universal_master_0_agent:rp_ready -> rsp_xbar_mux_002:src_ready
	wire          limiter_002_cmd_src_endofpacket;                                                                              // limiter_002:cmd_src_endofpacket -> cmd_xbar_demux_003:sink_endofpacket
	wire          limiter_002_cmd_src_startofpacket;                                                                            // limiter_002:cmd_src_startofpacket -> cmd_xbar_demux_003:sink_startofpacket
	wire  [112:0] limiter_002_cmd_src_data;                                                                                     // limiter_002:cmd_src_data -> cmd_xbar_demux_003:sink_data
	wire   [11:0] limiter_002_cmd_src_channel;                                                                                  // limiter_002:cmd_src_channel -> cmd_xbar_demux_003:sink_channel
	wire          limiter_002_cmd_src_ready;                                                                                    // cmd_xbar_demux_003:sink_ready -> limiter_002:cmd_src_ready
	wire          rsp_xbar_mux_003_src_endofpacket;                                                                             // rsp_xbar_mux_003:src_endofpacket -> limiter_002:rsp_sink_endofpacket
	wire          rsp_xbar_mux_003_src_valid;                                                                                   // rsp_xbar_mux_003:src_valid -> limiter_002:rsp_sink_valid
	wire          rsp_xbar_mux_003_src_startofpacket;                                                                           // rsp_xbar_mux_003:src_startofpacket -> limiter_002:rsp_sink_startofpacket
	wire  [112:0] rsp_xbar_mux_003_src_data;                                                                                    // rsp_xbar_mux_003:src_data -> limiter_002:rsp_sink_data
	wire   [11:0] rsp_xbar_mux_003_src_channel;                                                                                 // rsp_xbar_mux_003:src_channel -> limiter_002:rsp_sink_channel
	wire          rsp_xbar_mux_003_src_ready;                                                                                   // limiter_002:rsp_sink_ready -> rsp_xbar_mux_003:src_ready
	wire          addr_router_004_src_endofpacket;                                                                              // addr_router_004:src_endofpacket -> cmd_xbar_demux_004:sink_endofpacket
	wire          addr_router_004_src_valid;                                                                                    // addr_router_004:src_valid -> cmd_xbar_demux_004:sink_valid
	wire          addr_router_004_src_startofpacket;                                                                            // addr_router_004:src_startofpacket -> cmd_xbar_demux_004:sink_startofpacket
	wire  [112:0] addr_router_004_src_data;                                                                                     // addr_router_004:src_data -> cmd_xbar_demux_004:sink_data
	wire   [11:0] addr_router_004_src_channel;                                                                                  // addr_router_004:src_channel -> cmd_xbar_demux_004:sink_channel
	wire          addr_router_004_src_ready;                                                                                    // cmd_xbar_demux_004:sink_ready -> addr_router_004:src_ready
	wire          rsp_xbar_demux_001_src2_ready;                                                                                // ethernet_subsystem_sgdma_rx_m_write_translator_avalon_universal_master_0_agent:rp_ready -> rsp_xbar_demux_001:src2_ready
	wire          addr_router_005_src_endofpacket;                                                                              // addr_router_005:src_endofpacket -> cmd_xbar_demux_005:sink_endofpacket
	wire          addr_router_005_src_valid;                                                                                    // addr_router_005:src_valid -> cmd_xbar_demux_005:sink_valid
	wire          addr_router_005_src_startofpacket;                                                                            // addr_router_005:src_startofpacket -> cmd_xbar_demux_005:sink_startofpacket
	wire  [112:0] addr_router_005_src_data;                                                                                     // addr_router_005:src_data -> cmd_xbar_demux_005:sink_data
	wire   [11:0] addr_router_005_src_channel;                                                                                  // addr_router_005:src_channel -> cmd_xbar_demux_005:sink_channel
	wire          addr_router_005_src_ready;                                                                                    // cmd_xbar_demux_005:sink_ready -> addr_router_005:src_ready
	wire          rsp_xbar_demux_001_src3_ready;                                                                                // ethernet_subsystem_sgdma_tx_m_read_translator_avalon_universal_master_0_agent:rp_ready -> rsp_xbar_demux_001:src3_ready
	wire          cmd_xbar_mux_src_endofpacket;                                                                                 // cmd_xbar_mux:src_endofpacket -> burst_adapter:sink0_endofpacket
	wire          cmd_xbar_mux_src_valid;                                                                                       // cmd_xbar_mux:src_valid -> burst_adapter:sink0_valid
	wire          cmd_xbar_mux_src_startofpacket;                                                                               // cmd_xbar_mux:src_startofpacket -> burst_adapter:sink0_startofpacket
	wire  [112:0] cmd_xbar_mux_src_data;                                                                                        // cmd_xbar_mux:src_data -> burst_adapter:sink0_data
	wire   [11:0] cmd_xbar_mux_src_channel;                                                                                     // cmd_xbar_mux:src_channel -> burst_adapter:sink0_channel
	wire          cmd_xbar_mux_src_ready;                                                                                       // burst_adapter:sink0_ready -> cmd_xbar_mux:src_ready
	wire          id_router_src_endofpacket;                                                                                    // id_router:src_endofpacket -> rsp_xbar_demux:sink_endofpacket
	wire          id_router_src_valid;                                                                                          // id_router:src_valid -> rsp_xbar_demux:sink_valid
	wire          id_router_src_startofpacket;                                                                                  // id_router:src_startofpacket -> rsp_xbar_demux:sink_startofpacket
	wire  [112:0] id_router_src_data;                                                                                           // id_router:src_data -> rsp_xbar_demux:sink_data
	wire   [11:0] id_router_src_channel;                                                                                        // id_router:src_channel -> rsp_xbar_demux:sink_channel
	wire          id_router_src_ready;                                                                                          // rsp_xbar_demux:sink_ready -> id_router:src_ready
	wire          cmd_xbar_mux_001_src_endofpacket;                                                                             // cmd_xbar_mux_001:src_endofpacket -> burst_adapter_001:sink0_endofpacket
	wire          cmd_xbar_mux_001_src_valid;                                                                                   // cmd_xbar_mux_001:src_valid -> burst_adapter_001:sink0_valid
	wire          cmd_xbar_mux_001_src_startofpacket;                                                                           // cmd_xbar_mux_001:src_startofpacket -> burst_adapter_001:sink0_startofpacket
	wire  [112:0] cmd_xbar_mux_001_src_data;                                                                                    // cmd_xbar_mux_001:src_data -> burst_adapter_001:sink0_data
	wire   [11:0] cmd_xbar_mux_001_src_channel;                                                                                 // cmd_xbar_mux_001:src_channel -> burst_adapter_001:sink0_channel
	wire          cmd_xbar_mux_001_src_ready;                                                                                   // burst_adapter_001:sink0_ready -> cmd_xbar_mux_001:src_ready
	wire          id_router_001_src_endofpacket;                                                                                // id_router_001:src_endofpacket -> rsp_xbar_demux_001:sink_endofpacket
	wire          id_router_001_src_valid;                                                                                      // id_router_001:src_valid -> rsp_xbar_demux_001:sink_valid
	wire          id_router_001_src_startofpacket;                                                                              // id_router_001:src_startofpacket -> rsp_xbar_demux_001:sink_startofpacket
	wire  [112:0] id_router_001_src_data;                                                                                       // id_router_001:src_data -> rsp_xbar_demux_001:sink_data
	wire   [11:0] id_router_001_src_channel;                                                                                    // id_router_001:src_channel -> rsp_xbar_demux_001:sink_channel
	wire          id_router_001_src_ready;                                                                                      // rsp_xbar_demux_001:sink_ready -> id_router_001:src_ready
	wire          cmd_xbar_demux_001_src2_ready;                                                                                // burst_adapter_002:sink0_ready -> cmd_xbar_demux_001:src2_ready
	wire          id_router_002_src_endofpacket;                                                                                // id_router_002:src_endofpacket -> rsp_xbar_demux_002:sink_endofpacket
	wire          id_router_002_src_valid;                                                                                      // id_router_002:src_valid -> rsp_xbar_demux_002:sink_valid
	wire          id_router_002_src_startofpacket;                                                                              // id_router_002:src_startofpacket -> rsp_xbar_demux_002:sink_startofpacket
	wire  [112:0] id_router_002_src_data;                                                                                       // id_router_002:src_data -> rsp_xbar_demux_002:sink_data
	wire   [11:0] id_router_002_src_channel;                                                                                    // id_router_002:src_channel -> rsp_xbar_demux_002:sink_channel
	wire          id_router_002_src_ready;                                                                                      // rsp_xbar_demux_002:sink_ready -> id_router_002:src_ready
	wire          cmd_xbar_mux_003_src_endofpacket;                                                                             // cmd_xbar_mux_003:src_endofpacket -> burst_adapter_003:sink0_endofpacket
	wire          cmd_xbar_mux_003_src_valid;                                                                                   // cmd_xbar_mux_003:src_valid -> burst_adapter_003:sink0_valid
	wire          cmd_xbar_mux_003_src_startofpacket;                                                                           // cmd_xbar_mux_003:src_startofpacket -> burst_adapter_003:sink0_startofpacket
	wire  [112:0] cmd_xbar_mux_003_src_data;                                                                                    // cmd_xbar_mux_003:src_data -> burst_adapter_003:sink0_data
	wire   [11:0] cmd_xbar_mux_003_src_channel;                                                                                 // cmd_xbar_mux_003:src_channel -> burst_adapter_003:sink0_channel
	wire          cmd_xbar_mux_003_src_ready;                                                                                   // burst_adapter_003:sink0_ready -> cmd_xbar_mux_003:src_ready
	wire          id_router_003_src_endofpacket;                                                                                // id_router_003:src_endofpacket -> rsp_xbar_demux_003:sink_endofpacket
	wire          id_router_003_src_valid;                                                                                      // id_router_003:src_valid -> rsp_xbar_demux_003:sink_valid
	wire          id_router_003_src_startofpacket;                                                                              // id_router_003:src_startofpacket -> rsp_xbar_demux_003:sink_startofpacket
	wire  [112:0] id_router_003_src_data;                                                                                       // id_router_003:src_data -> rsp_xbar_demux_003:sink_data
	wire   [11:0] id_router_003_src_channel;                                                                                    // id_router_003:src_channel -> rsp_xbar_demux_003:sink_channel
	wire          id_router_003_src_ready;                                                                                      // rsp_xbar_demux_003:sink_ready -> id_router_003:src_ready
	wire          cmd_xbar_demux_001_src4_ready;                                                                                // burst_adapter_004:sink0_ready -> cmd_xbar_demux_001:src4_ready
	wire          id_router_004_src_endofpacket;                                                                                // id_router_004:src_endofpacket -> rsp_xbar_demux_004:sink_endofpacket
	wire          id_router_004_src_valid;                                                                                      // id_router_004:src_valid -> rsp_xbar_demux_004:sink_valid
	wire          id_router_004_src_startofpacket;                                                                              // id_router_004:src_startofpacket -> rsp_xbar_demux_004:sink_startofpacket
	wire  [112:0] id_router_004_src_data;                                                                                       // id_router_004:src_data -> rsp_xbar_demux_004:sink_data
	wire   [11:0] id_router_004_src_channel;                                                                                    // id_router_004:src_channel -> rsp_xbar_demux_004:sink_channel
	wire          id_router_004_src_ready;                                                                                      // rsp_xbar_demux_004:sink_ready -> id_router_004:src_ready
	wire          cmd_xbar_demux_001_src5_ready;                                                                                // burst_adapter_005:sink0_ready -> cmd_xbar_demux_001:src5_ready
	wire          id_router_005_src_endofpacket;                                                                                // id_router_005:src_endofpacket -> rsp_xbar_demux_005:sink_endofpacket
	wire          id_router_005_src_valid;                                                                                      // id_router_005:src_valid -> rsp_xbar_demux_005:sink_valid
	wire          id_router_005_src_startofpacket;                                                                              // id_router_005:src_startofpacket -> rsp_xbar_demux_005:sink_startofpacket
	wire  [112:0] id_router_005_src_data;                                                                                       // id_router_005:src_data -> rsp_xbar_demux_005:sink_data
	wire   [11:0] id_router_005_src_channel;                                                                                    // id_router_005:src_channel -> rsp_xbar_demux_005:sink_channel
	wire          id_router_005_src_ready;                                                                                      // rsp_xbar_demux_005:sink_ready -> id_router_005:src_ready
	wire          cmd_xbar_demux_001_src6_ready;                                                                                // burst_adapter_006:sink0_ready -> cmd_xbar_demux_001:src6_ready
	wire          id_router_006_src_endofpacket;                                                                                // id_router_006:src_endofpacket -> rsp_xbar_demux_006:sink_endofpacket
	wire          id_router_006_src_valid;                                                                                      // id_router_006:src_valid -> rsp_xbar_demux_006:sink_valid
	wire          id_router_006_src_startofpacket;                                                                              // id_router_006:src_startofpacket -> rsp_xbar_demux_006:sink_startofpacket
	wire  [112:0] id_router_006_src_data;                                                                                       // id_router_006:src_data -> rsp_xbar_demux_006:sink_data
	wire   [11:0] id_router_006_src_channel;                                                                                    // id_router_006:src_channel -> rsp_xbar_demux_006:sink_channel
	wire          id_router_006_src_ready;                                                                                      // rsp_xbar_demux_006:sink_ready -> id_router_006:src_ready
	wire          cmd_xbar_demux_001_src7_ready;                                                                                // burst_adapter_007:sink0_ready -> cmd_xbar_demux_001:src7_ready
	wire          id_router_007_src_endofpacket;                                                                                // id_router_007:src_endofpacket -> rsp_xbar_demux_007:sink_endofpacket
	wire          id_router_007_src_valid;                                                                                      // id_router_007:src_valid -> rsp_xbar_demux_007:sink_valid
	wire          id_router_007_src_startofpacket;                                                                              // id_router_007:src_startofpacket -> rsp_xbar_demux_007:sink_startofpacket
	wire  [112:0] id_router_007_src_data;                                                                                       // id_router_007:src_data -> rsp_xbar_demux_007:sink_data
	wire   [11:0] id_router_007_src_channel;                                                                                    // id_router_007:src_channel -> rsp_xbar_demux_007:sink_channel
	wire          id_router_007_src_ready;                                                                                      // rsp_xbar_demux_007:sink_ready -> id_router_007:src_ready
	wire          cmd_xbar_mux_008_src_endofpacket;                                                                             // cmd_xbar_mux_008:src_endofpacket -> carControl_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_mux_008_src_valid;                                                                                   // cmd_xbar_mux_008:src_valid -> carControl_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_mux_008_src_startofpacket;                                                                           // cmd_xbar_mux_008:src_startofpacket -> carControl_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [112:0] cmd_xbar_mux_008_src_data;                                                                                    // cmd_xbar_mux_008:src_data -> carControl_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_data
	wire   [11:0] cmd_xbar_mux_008_src_channel;                                                                                 // cmd_xbar_mux_008:src_channel -> carControl_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_mux_008_src_ready;                                                                                   // carControl_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_008:src_ready
	wire          id_router_008_src_endofpacket;                                                                                // id_router_008:src_endofpacket -> rsp_xbar_demux_008:sink_endofpacket
	wire          id_router_008_src_valid;                                                                                      // id_router_008:src_valid -> rsp_xbar_demux_008:sink_valid
	wire          id_router_008_src_startofpacket;                                                                              // id_router_008:src_startofpacket -> rsp_xbar_demux_008:sink_startofpacket
	wire  [112:0] id_router_008_src_data;                                                                                       // id_router_008:src_data -> rsp_xbar_demux_008:sink_data
	wire   [11:0] id_router_008_src_channel;                                                                                    // id_router_008:src_channel -> rsp_xbar_demux_008:sink_channel
	wire          id_router_008_src_ready;                                                                                      // rsp_xbar_demux_008:sink_ready -> id_router_008:src_ready
	wire          cmd_xbar_mux_009_src_endofpacket;                                                                             // cmd_xbar_mux_009:src_endofpacket -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_mux_009_src_valid;                                                                                   // cmd_xbar_mux_009:src_valid -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_mux_009_src_startofpacket;                                                                           // cmd_xbar_mux_009:src_startofpacket -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [112:0] cmd_xbar_mux_009_src_data;                                                                                    // cmd_xbar_mux_009:src_data -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [11:0] cmd_xbar_mux_009_src_channel;                                                                                 // cmd_xbar_mux_009:src_channel -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_mux_009_src_ready;                                                                                   // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_009:src_ready
	wire          id_router_009_src_endofpacket;                                                                                // id_router_009:src_endofpacket -> rsp_xbar_demux_009:sink_endofpacket
	wire          id_router_009_src_valid;                                                                                      // id_router_009:src_valid -> rsp_xbar_demux_009:sink_valid
	wire          id_router_009_src_startofpacket;                                                                              // id_router_009:src_startofpacket -> rsp_xbar_demux_009:sink_startofpacket
	wire  [112:0] id_router_009_src_data;                                                                                       // id_router_009:src_data -> rsp_xbar_demux_009:sink_data
	wire   [11:0] id_router_009_src_channel;                                                                                    // id_router_009:src_channel -> rsp_xbar_demux_009:sink_channel
	wire          id_router_009_src_ready;                                                                                      // rsp_xbar_demux_009:sink_ready -> id_router_009:src_ready
	wire          cmd_xbar_demux_002_src3_ready;                                                                                // jtaguart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_002:src3_ready
	wire          id_router_010_src_endofpacket;                                                                                // id_router_010:src_endofpacket -> rsp_xbar_demux_010:sink_endofpacket
	wire          id_router_010_src_valid;                                                                                      // id_router_010:src_valid -> rsp_xbar_demux_010:sink_valid
	wire          id_router_010_src_startofpacket;                                                                              // id_router_010:src_startofpacket -> rsp_xbar_demux_010:sink_startofpacket
	wire  [112:0] id_router_010_src_data;                                                                                       // id_router_010:src_data -> rsp_xbar_demux_010:sink_data
	wire   [11:0] id_router_010_src_channel;                                                                                    // id_router_010:src_channel -> rsp_xbar_demux_010:sink_channel
	wire          id_router_010_src_ready;                                                                                      // rsp_xbar_demux_010:sink_ready -> id_router_010:src_ready
	wire          cmd_xbar_demux_002_src4_ready;                                                                                // prio_arbiter_0_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_002:src4_ready
	wire          id_router_011_src_endofpacket;                                                                                // id_router_011:src_endofpacket -> rsp_xbar_demux_011:sink_endofpacket
	wire          id_router_011_src_valid;                                                                                      // id_router_011:src_valid -> rsp_xbar_demux_011:sink_valid
	wire          id_router_011_src_startofpacket;                                                                              // id_router_011:src_startofpacket -> rsp_xbar_demux_011:sink_startofpacket
	wire  [112:0] id_router_011_src_data;                                                                                       // id_router_011:src_data -> rsp_xbar_demux_011:sink_data
	wire   [11:0] id_router_011_src_channel;                                                                                    // id_router_011:src_channel -> rsp_xbar_demux_011:sink_channel
	wire          id_router_011_src_ready;                                                                                      // rsp_xbar_demux_011:sink_ready -> id_router_011:src_ready
	wire          cmd_xbar_demux_006_src0_endofpacket;                                                                          // cmd_xbar_demux_006:src0_endofpacket -> burst_adapter_008:sink0_endofpacket
	wire          cmd_xbar_demux_006_src0_valid;                                                                                // cmd_xbar_demux_006:src0_valid -> burst_adapter_008:sink0_valid
	wire          cmd_xbar_demux_006_src0_startofpacket;                                                                        // cmd_xbar_demux_006:src0_startofpacket -> burst_adapter_008:sink0_startofpacket
	wire  [102:0] cmd_xbar_demux_006_src0_data;                                                                                 // cmd_xbar_demux_006:src0_data -> burst_adapter_008:sink0_data
	wire    [0:0] cmd_xbar_demux_006_src0_channel;                                                                              // cmd_xbar_demux_006:src0_channel -> burst_adapter_008:sink0_channel
	wire          rsp_xbar_demux_012_src0_endofpacket;                                                                          // rsp_xbar_demux_012:src0_endofpacket -> traffic_gen_0_avalon_master_0_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire          rsp_xbar_demux_012_src0_valid;                                                                                // rsp_xbar_demux_012:src0_valid -> traffic_gen_0_avalon_master_0_translator_avalon_universal_master_0_agent:rp_valid
	wire          rsp_xbar_demux_012_src0_startofpacket;                                                                        // rsp_xbar_demux_012:src0_startofpacket -> traffic_gen_0_avalon_master_0_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [102:0] rsp_xbar_demux_012_src0_data;                                                                                 // rsp_xbar_demux_012:src0_data -> traffic_gen_0_avalon_master_0_translator_avalon_universal_master_0_agent:rp_data
	wire    [0:0] rsp_xbar_demux_012_src0_channel;                                                                              // rsp_xbar_demux_012:src0_channel -> traffic_gen_0_avalon_master_0_translator_avalon_universal_master_0_agent:rp_channel
	wire          addr_router_006_src_endofpacket;                                                                              // addr_router_006:src_endofpacket -> cmd_xbar_demux_006:sink_endofpacket
	wire          addr_router_006_src_valid;                                                                                    // addr_router_006:src_valid -> cmd_xbar_demux_006:sink_valid
	wire          addr_router_006_src_startofpacket;                                                                            // addr_router_006:src_startofpacket -> cmd_xbar_demux_006:sink_startofpacket
	wire  [102:0] addr_router_006_src_data;                                                                                     // addr_router_006:src_data -> cmd_xbar_demux_006:sink_data
	wire    [0:0] addr_router_006_src_channel;                                                                                  // addr_router_006:src_channel -> cmd_xbar_demux_006:sink_channel
	wire          addr_router_006_src_ready;                                                                                    // cmd_xbar_demux_006:sink_ready -> addr_router_006:src_ready
	wire          rsp_xbar_demux_012_src0_ready;                                                                                // traffic_gen_0_avalon_master_0_translator_avalon_universal_master_0_agent:rp_ready -> rsp_xbar_demux_012:src0_ready
	wire          cmd_xbar_demux_006_src0_ready;                                                                                // burst_adapter_008:sink0_ready -> cmd_xbar_demux_006:src0_ready
	wire          id_router_012_src_endofpacket;                                                                                // id_router_012:src_endofpacket -> rsp_xbar_demux_012:sink_endofpacket
	wire          id_router_012_src_valid;                                                                                      // id_router_012:src_valid -> rsp_xbar_demux_012:sink_valid
	wire          id_router_012_src_startofpacket;                                                                              // id_router_012:src_startofpacket -> rsp_xbar_demux_012:sink_startofpacket
	wire  [102:0] id_router_012_src_data;                                                                                       // id_router_012:src_data -> rsp_xbar_demux_012:sink_data
	wire    [0:0] id_router_012_src_channel;                                                                                    // id_router_012:src_channel -> rsp_xbar_demux_012:sink_channel
	wire          id_router_012_src_ready;                                                                                      // rsp_xbar_demux_012:sink_ready -> id_router_012:src_ready
	wire          cmd_xbar_demux_007_src0_endofpacket;                                                                          // cmd_xbar_demux_007:src0_endofpacket -> burst_adapter_009:sink0_endofpacket
	wire          cmd_xbar_demux_007_src0_valid;                                                                                // cmd_xbar_demux_007:src0_valid -> burst_adapter_009:sink0_valid
	wire          cmd_xbar_demux_007_src0_startofpacket;                                                                        // cmd_xbar_demux_007:src0_startofpacket -> burst_adapter_009:sink0_startofpacket
	wire  [102:0] cmd_xbar_demux_007_src0_data;                                                                                 // cmd_xbar_demux_007:src0_data -> burst_adapter_009:sink0_data
	wire    [0:0] cmd_xbar_demux_007_src0_channel;                                                                              // cmd_xbar_demux_007:src0_channel -> burst_adapter_009:sink0_channel
	wire          rsp_xbar_demux_013_src0_endofpacket;                                                                          // rsp_xbar_demux_013:src0_endofpacket -> traffic_gen_1_avalon_master_0_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire          rsp_xbar_demux_013_src0_valid;                                                                                // rsp_xbar_demux_013:src0_valid -> traffic_gen_1_avalon_master_0_translator_avalon_universal_master_0_agent:rp_valid
	wire          rsp_xbar_demux_013_src0_startofpacket;                                                                        // rsp_xbar_demux_013:src0_startofpacket -> traffic_gen_1_avalon_master_0_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [102:0] rsp_xbar_demux_013_src0_data;                                                                                 // rsp_xbar_demux_013:src0_data -> traffic_gen_1_avalon_master_0_translator_avalon_universal_master_0_agent:rp_data
	wire    [0:0] rsp_xbar_demux_013_src0_channel;                                                                              // rsp_xbar_demux_013:src0_channel -> traffic_gen_1_avalon_master_0_translator_avalon_universal_master_0_agent:rp_channel
	wire          addr_router_007_src_endofpacket;                                                                              // addr_router_007:src_endofpacket -> cmd_xbar_demux_007:sink_endofpacket
	wire          addr_router_007_src_valid;                                                                                    // addr_router_007:src_valid -> cmd_xbar_demux_007:sink_valid
	wire          addr_router_007_src_startofpacket;                                                                            // addr_router_007:src_startofpacket -> cmd_xbar_demux_007:sink_startofpacket
	wire  [102:0] addr_router_007_src_data;                                                                                     // addr_router_007:src_data -> cmd_xbar_demux_007:sink_data
	wire    [0:0] addr_router_007_src_channel;                                                                                  // addr_router_007:src_channel -> cmd_xbar_demux_007:sink_channel
	wire          addr_router_007_src_ready;                                                                                    // cmd_xbar_demux_007:sink_ready -> addr_router_007:src_ready
	wire          rsp_xbar_demux_013_src0_ready;                                                                                // traffic_gen_1_avalon_master_0_translator_avalon_universal_master_0_agent:rp_ready -> rsp_xbar_demux_013:src0_ready
	wire          cmd_xbar_demux_007_src0_ready;                                                                                // burst_adapter_009:sink0_ready -> cmd_xbar_demux_007:src0_ready
	wire          id_router_013_src_endofpacket;                                                                                // id_router_013:src_endofpacket -> rsp_xbar_demux_013:sink_endofpacket
	wire          id_router_013_src_valid;                                                                                      // id_router_013:src_valid -> rsp_xbar_demux_013:sink_valid
	wire          id_router_013_src_startofpacket;                                                                              // id_router_013:src_startofpacket -> rsp_xbar_demux_013:sink_startofpacket
	wire  [102:0] id_router_013_src_data;                                                                                       // id_router_013:src_data -> rsp_xbar_demux_013:sink_data
	wire    [0:0] id_router_013_src_channel;                                                                                    // id_router_013:src_channel -> rsp_xbar_demux_013:sink_channel
	wire          id_router_013_src_ready;                                                                                      // rsp_xbar_demux_013:sink_ready -> id_router_013:src_ready
	wire   [11:0] limiter_cmd_valid_data;                                                                                       // limiter:cmd_src_valid -> cmd_xbar_demux:sink_valid
	wire   [11:0] limiter_001_cmd_valid_data;                                                                                   // limiter_001:cmd_src_valid -> cmd_xbar_demux_001:sink_valid
	wire   [11:0] limiter_002_cmd_valid_data;                                                                                   // limiter_002:cmd_src_valid -> cmd_xbar_demux_003:sink_valid
	wire          irq_mapper_receiver0_irq;                                                                                     // jtaguart_0:av_irq -> irq_mapper:receiver0_irq
	wire          irq_mapper_receiver1_irq;                                                                                     // com_timer:irq -> irq_mapper:receiver1_irq
	wire          irq_mapper_receiver2_irq;                                                                                     // ethernet_subsystem:sgdma_rx_csr_irq_irq -> irq_mapper:receiver2_irq
	wire          irq_mapper_receiver3_irq;                                                                                     // ethernet_subsystem:sgdma_tx_csr_irq_irq -> irq_mapper:receiver3_irq
	wire   [31:0] com_nios_d_irq_irq;                                                                                           // irq_mapper:sender_irq -> com_nios:d_irq
	wire          irq_mapper_001_receiver0_irq;                                                                                 // jtaguart_1:av_irq -> irq_mapper_001:receiver0_irq
	wire   [31:0] carcontrol_nios_d_irq_irq;                                                                                    // irq_mapper_001:sender_irq -> carControl_nios:d_irq

	nios_system_com_nios com_nios (
		.clk                                   (clk_clk),                                                                 //                       clk.clk
		.reset_n                               (~rst_controller_reset_out_reset),                                         //                   reset_n.reset_n
		.d_address                             (com_nios_data_master_address),                                            //               data_master.address
		.d_byteenable                          (com_nios_data_master_byteenable),                                         //                          .byteenable
		.d_read                                (com_nios_data_master_read),                                               //                          .read
		.d_readdata                            (com_nios_data_master_readdata),                                           //                          .readdata
		.d_waitrequest                         (com_nios_data_master_waitrequest),                                        //                          .waitrequest
		.d_write                               (com_nios_data_master_write),                                              //                          .write
		.d_writedata                           (com_nios_data_master_writedata),                                          //                          .writedata
		.d_burstcount                          (com_nios_data_master_burstcount),                                         //                          .burstcount
		.d_readdatavalid                       (com_nios_data_master_readdatavalid),                                      //                          .readdatavalid
		.jtag_debug_module_debugaccess_to_roms (com_nios_data_master_debugaccess),                                        //                          .debugaccess
		.i_address                             (com_nios_instruction_master_address),                                     //        instruction_master.address
		.i_read                                (com_nios_instruction_master_read),                                        //                          .read
		.i_readdata                            (com_nios_instruction_master_readdata),                                    //                          .readdata
		.i_waitrequest                         (com_nios_instruction_master_waitrequest),                                 //                          .waitrequest
		.i_burstcount                          (com_nios_instruction_master_burstcount),                                  //                          .burstcount
		.i_readdatavalid                       (com_nios_instruction_master_readdatavalid),                               //                          .readdatavalid
		.d_irq                                 (com_nios_d_irq_irq),                                                      //                     d_irq.irq
		.jtag_debug_module_resetrequest        (com_nios_jtag_debug_module_reset_reset),                                  //   jtag_debug_module_reset.reset
		.jtag_debug_module_address             (com_nios_jtag_debug_module_translator_avalon_anti_slave_0_address),       //         jtag_debug_module.address
		.jtag_debug_module_begintransfer       (com_nios_jtag_debug_module_translator_avalon_anti_slave_0_begintransfer), //                          .begintransfer
		.jtag_debug_module_byteenable          (com_nios_jtag_debug_module_translator_avalon_anti_slave_0_byteenable),    //                          .byteenable
		.jtag_debug_module_debugaccess         (com_nios_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess),   //                          .debugaccess
		.jtag_debug_module_readdata            (com_nios_jtag_debug_module_translator_avalon_anti_slave_0_readdata),      //                          .readdata
		.jtag_debug_module_select              (com_nios_jtag_debug_module_translator_avalon_anti_slave_0_chipselect),    //                          .chipselect
		.jtag_debug_module_write               (com_nios_jtag_debug_module_translator_avalon_anti_slave_0_write),         //                          .write
		.jtag_debug_module_writedata           (com_nios_jtag_debug_module_translator_avalon_anti_slave_0_writedata),     //                          .writedata
		.no_ci_readra                          ()                                                                         // custom_instruction_master.readra
	);

	nios_system_jtaguart_0 jtaguart_0 (
		.clk            (clk_clk),                                                                 //               clk.clk
		.rst_n          (~rst_controller_001_reset_out_reset),                                     //             reset.reset_n
		.av_chipselect  (jtaguart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (jtaguart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_address),     //                  .address
		.av_read_n      (~jtaguart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_read),       //                  .read_n
		.av_readdata    (jtaguart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata),    //                  .readdata
		.av_write_n     (~jtaguart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_write),      //                  .write_n
		.av_writedata   (jtaguart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata),   //                  .writedata
		.av_waitrequest (jtaguart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                                                 //               irq.irq
	);

	nios_system_carControl_nios carcontrol_nios (
		.clk                                   (clk_clk),                                                                        //                       clk.clk
		.reset_n                               (~rst_controller_reset_out_reset),                                                //                   reset_n.reset_n
		.d_address                             (carcontrol_nios_data_master_address),                                            //               data_master.address
		.d_byteenable                          (carcontrol_nios_data_master_byteenable),                                         //                          .byteenable
		.d_read                                (carcontrol_nios_data_master_read),                                               //                          .read
		.d_readdata                            (carcontrol_nios_data_master_readdata),                                           //                          .readdata
		.d_waitrequest                         (carcontrol_nios_data_master_waitrequest),                                        //                          .waitrequest
		.d_write                               (carcontrol_nios_data_master_write),                                              //                          .write
		.d_writedata                           (carcontrol_nios_data_master_writedata),                                          //                          .writedata
		.jtag_debug_module_debugaccess_to_roms (carcontrol_nios_data_master_debugaccess),                                        //                          .debugaccess
		.i_address                             (carcontrol_nios_instruction_master_address),                                     //        instruction_master.address
		.i_read                                (carcontrol_nios_instruction_master_read),                                        //                          .read
		.i_readdata                            (carcontrol_nios_instruction_master_readdata),                                    //                          .readdata
		.i_waitrequest                         (carcontrol_nios_instruction_master_waitrequest),                                 //                          .waitrequest
		.i_readdatavalid                       (carcontrol_nios_instruction_master_readdatavalid),                               //                          .readdatavalid
		.d_irq                                 (carcontrol_nios_d_irq_irq),                                                      //                     d_irq.irq
		.jtag_debug_module_resetrequest        (carcontrol_nios_jtag_debug_module_reset_reset),                                  //   jtag_debug_module_reset.reset
		.jtag_debug_module_address             (carcontrol_nios_jtag_debug_module_translator_avalon_anti_slave_0_address),       //         jtag_debug_module.address
		.jtag_debug_module_begintransfer       (carcontrol_nios_jtag_debug_module_translator_avalon_anti_slave_0_begintransfer), //                          .begintransfer
		.jtag_debug_module_byteenable          (carcontrol_nios_jtag_debug_module_translator_avalon_anti_slave_0_byteenable),    //                          .byteenable
		.jtag_debug_module_debugaccess         (carcontrol_nios_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess),   //                          .debugaccess
		.jtag_debug_module_readdata            (carcontrol_nios_jtag_debug_module_translator_avalon_anti_slave_0_readdata),      //                          .readdata
		.jtag_debug_module_select              (carcontrol_nios_jtag_debug_module_translator_avalon_anti_slave_0_chipselect),    //                          .chipselect
		.jtag_debug_module_write               (carcontrol_nios_jtag_debug_module_translator_avalon_anti_slave_0_write),         //                          .write
		.jtag_debug_module_writedata           (carcontrol_nios_jtag_debug_module_translator_avalon_anti_slave_0_writedata),     //                          .writedata
		.no_ci_readra                          ()                                                                                // custom_instruction_master.readra
	);

	nios_system_shared_memory shared_memory (
		.clk        (clk_clk),                                                    //   clk1.clk
		.address    (shared_memory_s1_translator_avalon_anti_slave_0_address),    //     s1.address
		.chipselect (shared_memory_s1_translator_avalon_anti_slave_0_chipselect), //       .chipselect
		.clken      (shared_memory_s1_translator_avalon_anti_slave_0_clken),      //       .clken
		.readdata   (shared_memory_s1_translator_avalon_anti_slave_0_readdata),   //       .readdata
		.write      (shared_memory_s1_translator_avalon_anti_slave_0_write),      //       .write
		.writedata  (shared_memory_s1_translator_avalon_anti_slave_0_writedata),  //       .writedata
		.byteenable (shared_memory_s1_translator_avalon_anti_slave_0_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset)                              // reset1.reset
	);

	nios_system_shared_memory_mutex shared_memory_mutex (
		.clk           (clk_clk),                                                          //   clk.clk
		.reset_n       (~rst_controller_reset_out_reset),                                  // reset.reset_n
		.address       (shared_memory_mutex_s1_translator_avalon_anti_slave_0_address),    //    s1.address
		.chipselect    (shared_memory_mutex_s1_translator_avalon_anti_slave_0_chipselect), //      .chipselect
		.data_from_cpu (shared_memory_mutex_s1_translator_avalon_anti_slave_0_writedata),  //      .writedata
		.data_to_cpu   (shared_memory_mutex_s1_translator_avalon_anti_slave_0_readdata),   //      .readdata
		.read          (shared_memory_mutex_s1_translator_avalon_anti_slave_0_read),       //      .read
		.write         (shared_memory_mutex_s1_translator_avalon_anti_slave_0_write)       //      .write
	);

	nios_system_com_timer com_timer (
		.clk        (clk_clk),                                                //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                        // reset.reset_n
		.address    (com_timer_s1_translator_avalon_anti_slave_0_address),    //    s1.address
		.writedata  (com_timer_s1_translator_avalon_anti_slave_0_writedata),  //      .writedata
		.readdata   (com_timer_s1_translator_avalon_anti_slave_0_readdata),   //      .readdata
		.chipselect (com_timer_s1_translator_avalon_anti_slave_0_chipselect), //      .chipselect
		.write_n    (~com_timer_s1_translator_avalon_anti_slave_0_write),     //      .write_n
		.irq        (irq_mapper_receiver1_irq)                                //   irq.irq
	);

	nios_system_com_memory com_memory (
		.clk            (clk_clk),                                                    //   clk.clk
		.reset_n        (~rst_controller_reset_out_reset),                            // reset.reset_n
		.az_addr        (com_memory_s1_translator_avalon_anti_slave_0_address),       //    s1.address
		.az_be_n        (~com_memory_s1_translator_avalon_anti_slave_0_byteenable),   //      .byteenable_n
		.az_cs          (com_memory_s1_translator_avalon_anti_slave_0_chipselect),    //      .chipselect
		.az_data        (com_memory_s1_translator_avalon_anti_slave_0_writedata),     //      .writedata
		.az_rd_n        (~com_memory_s1_translator_avalon_anti_slave_0_read),         //      .read_n
		.az_wr_n        (~com_memory_s1_translator_avalon_anti_slave_0_write),        //      .write_n
		.za_data        (com_memory_s1_translator_avalon_anti_slave_0_readdata),      //      .readdata
		.za_valid       (com_memory_s1_translator_avalon_anti_slave_0_readdatavalid), //      .readdatavalid
		.za_waitrequest (com_memory_s1_translator_avalon_anti_slave_0_waitrequest),   //      .waitrequest
		.zs_addr        (com_sdram_wire_addr),                                        //  wire.export
		.zs_ba          (com_sdram_wire_ba),                                          //      .export
		.zs_cas_n       (com_sdram_wire_cas_n),                                       //      .export
		.zs_cke         (com_sdram_wire_cke),                                         //      .export
		.zs_cs_n        (com_sdram_wire_cs_n),                                        //      .export
		.zs_dq          (com_sdram_wire_dq),                                          //      .export
		.zs_dqm         (com_sdram_wire_dqm),                                         //      .export
		.zs_ras_n       (com_sdram_wire_ras_n),                                       //      .export
		.zs_we_n        (com_sdram_wire_we_n)                                         //      .export
	);

	nios_system_onchip_memory2_0 onchip_memory2_0 (
		.clk        (clk_clk),                                                       //   clk1.clk
		.address    (onchip_memory2_0_s1_translator_avalon_anti_slave_0_address),    //     s1.address
		.chipselect (onchip_memory2_0_s1_translator_avalon_anti_slave_0_chipselect), //       .chipselect
		.clken      (onchip_memory2_0_s1_translator_avalon_anti_slave_0_clken),      //       .clken
		.readdata   (onchip_memory2_0_s1_translator_avalon_anti_slave_0_readdata),   //       .readdata
		.write      (onchip_memory2_0_s1_translator_avalon_anti_slave_0_write),      //       .write
		.writedata  (onchip_memory2_0_s1_translator_avalon_anti_slave_0_writedata),  //       .writedata
		.byteenable (onchip_memory2_0_s1_translator_avalon_anti_slave_0_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset)                                 // reset1.reset
	);

	nios_system_ethernet_subsystem ethernet_subsystem (
		.ethernet_subsys_clk_in_clk        (clk_clk),                                                                            //   ethernet_subsys_clk_in.clk
		.ethernet_subsys_reset_in_reset_n  (reset_reset_n),                                                                      // ethernet_subsys_reset_in.reset_n
		.ethernet_bridge_s0_waitrequest    (ethernet_subsystem_ethernet_bridge_s0_translator_avalon_anti_slave_0_waitrequest),   //       ethernet_bridge_s0.waitrequest
		.ethernet_bridge_s0_readdata       (ethernet_subsystem_ethernet_bridge_s0_translator_avalon_anti_slave_0_readdata),      //                         .readdata
		.ethernet_bridge_s0_readdatavalid  (ethernet_subsystem_ethernet_bridge_s0_translator_avalon_anti_slave_0_readdatavalid), //                         .readdatavalid
		.ethernet_bridge_s0_burstcount     (ethernet_subsystem_ethernet_bridge_s0_translator_avalon_anti_slave_0_burstcount),    //                         .burstcount
		.ethernet_bridge_s0_writedata      (ethernet_subsystem_ethernet_bridge_s0_translator_avalon_anti_slave_0_writedata),     //                         .writedata
		.ethernet_bridge_s0_address        (ethernet_subsystem_ethernet_bridge_s0_translator_avalon_anti_slave_0_address),       //                         .address
		.ethernet_bridge_s0_write          (ethernet_subsystem_ethernet_bridge_s0_translator_avalon_anti_slave_0_write),         //                         .write
		.ethernet_bridge_s0_read           (ethernet_subsystem_ethernet_bridge_s0_translator_avalon_anti_slave_0_read),          //                         .read
		.ethernet_bridge_s0_byteenable     (ethernet_subsystem_ethernet_bridge_s0_translator_avalon_anti_slave_0_byteenable),    //                         .byteenable
		.ethernet_bridge_s0_debugaccess    (ethernet_subsystem_ethernet_bridge_s0_translator_avalon_anti_slave_0_debugaccess),   //                         .debugaccess
		.tse_conduit_connection_rgmii_in   (tse_conduit_connection_rgmii_in),                                                    //   tse_conduit_connection.rgmii_in
		.tse_conduit_connection_rgmii_out  (tse_conduit_connection_rgmii_out),                                                   //                         .rgmii_out
		.tse_conduit_connection_rx_control (tse_conduit_connection_rx_control),                                                  //                         .rx_control
		.tse_conduit_connection_tx_control (tse_conduit_connection_tx_control),                                                  //                         .tx_control
		.tse_conduit_connection_tx_clk     (tse_conduit_connection_tx_clk),                                                      //                         .tx_clk
		.tse_conduit_connection_rx_clk     (tse_conduit_connection_rx_clk),                                                      //                         .rx_clk
		.tse_conduit_connection_set_10     (tse_conduit_connection_set_10),                                                      //                         .set_10
		.tse_conduit_connection_set_1000   (tse_conduit_connection_set_1000),                                                    //                         .set_1000
		.tse_conduit_connection_ena_10     (tse_conduit_connection_ena_10),                                                      //                         .ena_10
		.tse_conduit_connection_eth_mode   (tse_conduit_connection_eth_mode),                                                    //                         .eth_mode
		.tse_conduit_connection_mdio_out   (tse_conduit_connection_mdio_out),                                                    //                         .mdio_out
		.tse_conduit_connection_mdio_oen   (tse_conduit_connection_mdio_oen),                                                    //                         .mdio_oen
		.tse_conduit_connection_mdio_in    (tse_conduit_connection_mdio_in),                                                     //                         .mdio_in
		.tse_conduit_connection_mdc        (tse_conduit_connection_mdc),                                                         //                         .mdc
		.sgdma_rx_csr_irq_irq              (irq_mapper_receiver2_irq),                                                           //         sgdma_rx_csr_irq.irq
		.sgdma_rx_m_write_waitrequest      (ethernet_subsystem_sgdma_rx_m_write_waitrequest),                                    //         sgdma_rx_m_write.waitrequest
		.sgdma_rx_m_write_address          (ethernet_subsystem_sgdma_rx_m_write_address),                                        //                         .address
		.sgdma_rx_m_write_write            (ethernet_subsystem_sgdma_rx_m_write_write),                                          //                         .write
		.sgdma_rx_m_write_writedata        (ethernet_subsystem_sgdma_rx_m_write_writedata),                                      //                         .writedata
		.sgdma_rx_m_write_byteenable       (ethernet_subsystem_sgdma_rx_m_write_byteenable),                                     //                         .byteenable
		.sgdma_tx_csr_irq_irq              (irq_mapper_receiver3_irq),                                                           //         sgdma_tx_csr_irq.irq
		.sgdma_tx_m_read_readdata          (ethernet_subsystem_sgdma_tx_m_read_readdata),                                        //          sgdma_tx_m_read.readdata
		.sgdma_tx_m_read_readdatavalid     (ethernet_subsystem_sgdma_tx_m_read_readdatavalid),                                   //                         .readdatavalid
		.sgdma_tx_m_read_waitrequest       (ethernet_subsystem_sgdma_tx_m_read_waitrequest),                                     //                         .waitrequest
		.sgdma_tx_m_read_address           (ethernet_subsystem_sgdma_tx_m_read_address),                                         //                         .address
		.sgdma_tx_m_read_read              (ethernet_subsystem_sgdma_tx_m_read_read),                                            //                         .read
		.descriptor_memory_s2_address      (ethernet_subsystem_descriptor_memory_s2_translator_avalon_anti_slave_0_address),     //     descriptor_memory_s2.address
		.descriptor_memory_s2_chipselect   (ethernet_subsystem_descriptor_memory_s2_translator_avalon_anti_slave_0_chipselect),  //                         .chipselect
		.descriptor_memory_s2_clken        (ethernet_subsystem_descriptor_memory_s2_translator_avalon_anti_slave_0_clken),       //                         .clken
		.descriptor_memory_s2_readdata     (ethernet_subsystem_descriptor_memory_s2_translator_avalon_anti_slave_0_readdata),    //                         .readdata
		.descriptor_memory_s2_write        (ethernet_subsystem_descriptor_memory_s2_translator_avalon_anti_slave_0_write),       //                         .write
		.descriptor_memory_s2_writedata    (ethernet_subsystem_descriptor_memory_s2_translator_avalon_anti_slave_0_writedata),   //                         .writedata
		.descriptor_memory_s2_byteenable   (ethernet_subsystem_descriptor_memory_s2_translator_avalon_anti_slave_0_byteenable)   //                         .byteenable
	);

	nios_system_jtaguart_1 jtaguart_1 (
		.clk            (clk_clk),                                                                 //               clk.clk
		.rst_n          (~rst_controller_002_reset_out_reset),                                     //             reset.reset_n
		.av_chipselect  (jtaguart_1_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (jtaguart_1_avalon_jtag_slave_translator_avalon_anti_slave_0_address),     //                  .address
		.av_read_n      (~jtaguart_1_avalon_jtag_slave_translator_avalon_anti_slave_0_read),       //                  .read_n
		.av_readdata    (jtaguart_1_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata),    //                  .readdata
		.av_write_n     (~jtaguart_1_avalon_jtag_slave_translator_avalon_anti_slave_0_write),      //                  .write_n
		.av_writedata   (jtaguart_1_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata),   //                  .writedata
		.av_waitrequest (jtaguart_1_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_001_receiver0_irq)                                             //               irq.irq
	);

	prio_arbiter #(
		.SLAVE_ADDR_WIDTH     (26),
		.DATA_WIDTH           (32),
		.MASTER_ADDR_WIDTH    (28),
		.BYTE_ENABLE_BITS     (4),
		.NUM_OF_MASTERS       (4),
		.REQUEST_QUEUE_LENGTH (24),
		.SLOT_TIME            (1)
	) prio_arbiter_0 (
		.AVS_S0_CHIPSELECT      (prio_arbiter_0_s0_translator_avalon_anti_slave_0_chipselect),    //               s0.chipselect
		.AVS_S0_WRITE           (prio_arbiter_0_s0_translator_avalon_anti_slave_0_write),         //                 .write
		.AVS_S0_READ            (prio_arbiter_0_s0_translator_avalon_anti_slave_0_read),          //                 .read
		.AVS_S0_WRITEDATA       (prio_arbiter_0_s0_translator_avalon_anti_slave_0_writedata),     //                 .writedata
		.AVS_S0_BYTEENABLE      (prio_arbiter_0_s0_translator_avalon_anti_slave_0_byteenable),    //                 .byteenable
		.AVS_S0_READDATA        (prio_arbiter_0_s0_translator_avalon_anti_slave_0_readdata),      //                 .readdata
		.AVS_S0_READDATAVALID   (prio_arbiter_0_s0_translator_avalon_anti_slave_0_readdatavalid), //                 .readdatavalid
		.AVS_S0_WAITREQUEST     (prio_arbiter_0_s0_translator_avalon_anti_slave_0_waitrequest),   //                 .waitrequest
		.AVS_S0_ADDRESS         (prio_arbiter_0_s0_translator_avalon_anti_slave_0_address),       //                 .address
		.AVS_S1_ADDRESS         (prio_arbiter_0_s1_translator_avalon_anti_slave_0_address),       //               s1.address
		.AVS_S1_CHIPSELECT      (prio_arbiter_0_s1_translator_avalon_anti_slave_0_chipselect),    //                 .chipselect
		.AVS_S1_WRITE           (prio_arbiter_0_s1_translator_avalon_anti_slave_0_write),         //                 .write
		.AVS_S1_READ            (prio_arbiter_0_s1_translator_avalon_anti_slave_0_read),          //                 .read
		.AVS_S1_WRITEDATA       (prio_arbiter_0_s1_translator_avalon_anti_slave_0_writedata),     //                 .writedata
		.AVS_S1_BYTEENABLE      (prio_arbiter_0_s1_translator_avalon_anti_slave_0_byteenable),    //                 .byteenable
		.AVS_S1_READDATA        (prio_arbiter_0_s1_translator_avalon_anti_slave_0_readdata),      //                 .readdata
		.AVS_S1_READDATAVALID   (prio_arbiter_0_s1_translator_avalon_anti_slave_0_readdatavalid), //                 .readdatavalid
		.AVS_S1_WAITREQUEST     (prio_arbiter_0_s1_translator_avalon_anti_slave_0_waitrequest),   //                 .waitrequest
		.AVS_S2_ADDRESS         (prio_arbiter_0_s2_translator_avalon_anti_slave_0_address),       //               s2.address
		.AVS_S2_CHIPSELECT      (prio_arbiter_0_s2_translator_avalon_anti_slave_0_chipselect),    //                 .chipselect
		.AVS_S2_WRITE           (prio_arbiter_0_s2_translator_avalon_anti_slave_0_write),         //                 .write
		.AVS_S2_READ            (prio_arbiter_0_s2_translator_avalon_anti_slave_0_read),          //                 .read
		.AVS_S2_WRITEDATA       (prio_arbiter_0_s2_translator_avalon_anti_slave_0_writedata),     //                 .writedata
		.AVS_S2_BYTEENABLE      (prio_arbiter_0_s2_translator_avalon_anti_slave_0_byteenable),    //                 .byteenable
		.AVS_S2_READDATA        (prio_arbiter_0_s2_translator_avalon_anti_slave_0_readdata),      //                 .readdata
		.AVS_S2_READDATAVALID   (prio_arbiter_0_s2_translator_avalon_anti_slave_0_readdatavalid), //                 .readdatavalid
		.AVS_S2_WAITREQUEST     (prio_arbiter_0_s2_translator_avalon_anti_slave_0_waitrequest),   //                 .waitrequest
		.AVS_S3_ADDRESS         (prio_arbiter_0_s3_translator_avalon_anti_slave_0_address),       //               s3.address
		.AVS_S3_CHIPSELECT      (prio_arbiter_0_s3_translator_avalon_anti_slave_0_chipselect),    //                 .chipselect
		.AVS_S3_WRITE           (prio_arbiter_0_s3_translator_avalon_anti_slave_0_write),         //                 .write
		.AVS_S3_READ            (prio_arbiter_0_s3_translator_avalon_anti_slave_0_read),          //                 .read
		.AVS_S3_WRITEDATA       (prio_arbiter_0_s3_translator_avalon_anti_slave_0_writedata),     //                 .writedata
		.AVS_S3_BYTEENABLE      (prio_arbiter_0_s3_translator_avalon_anti_slave_0_byteenable),    //                 .byteenable
		.AVS_S3_READDATA        (prio_arbiter_0_s3_translator_avalon_anti_slave_0_readdata),      //                 .readdata
		.AVS_S3_READDATAVALID   (prio_arbiter_0_s3_translator_avalon_anti_slave_0_readdatavalid), //                 .readdatavalid
		.AVS_S3_WAITREQUEST     (prio_arbiter_0_s3_translator_avalon_anti_slave_0_waitrequest),   //                 .waitrequest
		.AVM_M1_ADDRESS         (prio_arbiter_0_m1_address),                                      //               m1.address
		.AVM_M1_READ            (prio_arbiter_0_m1_read),                                         //                 .read
		.AVM_M1_WRITE           (prio_arbiter_0_m1_write),                                        //                 .write
		.AVM_M1_WRITEDATA       (prio_arbiter_0_m1_writedata),                                    //                 .writedata
		.AVM_M1_BYTEENABLE      (prio_arbiter_0_m1_byteenable),                                   //                 .byteenable
		.AVM_M1_READDATA        (prio_arbiter_0_m1_readdata),                                     //                 .readdata
		.AVM_M1_WAITREQUEST     (prio_arbiter_0_m1_waitrequest),                                  //                 .waitrequest
		.AVM_M1_READDATAVALID   (prio_arbiter_0_m1_readdatavalid),                                //                 .readdatavalid
		.csi_clockreset_CLK     (clk_clk),                                                        //       clock_sink.clk
		.csi_clockreset_RESET_n (~rst_controller_reset_out_reset)                                 // clockreset_reset.reset_n
	);

	traffic_gen #(
		.SLAVE_ADDR_WIDTH  (26),
		.DATA_WIDTH        (32),
		.MASTER_ADDR_WIDTH (28),
		.BYTE_ENABLE_BITS  (4),
		.BURST_COUNT_BITS  (4),
		.BURST_LENGTH      (8),
		.NUM_OF_MASTERS    (4),
		.master_index      (1),
		.sopc_enable       (1)
	) traffic_gen_0 (
		.MASTER_ADDRES_AVM        (traffic_gen_0_avalon_master_0_address),       // avalon_master_0.address
		.MASTER_READ_AVM          (traffic_gen_0_avalon_master_0_read),          //                .read
		.MASTER_WRITE_AVM         (traffic_gen_0_avalon_master_0_write),         //                .write
		.MASTER_WRITEDATA_AVM     (traffic_gen_0_avalon_master_0_writedata),     //                .writedata
		.MASTER_BYTEENABLE_AVM    (traffic_gen_0_avalon_master_0_byteenable),    //                .byteenable
		.MASTER_READ_DATA_AVM     (traffic_gen_0_avalon_master_0_readdata),      //                .readdata
		.MASTER_WAITREQUEST_AVM   (traffic_gen_0_avalon_master_0_waitrequest),   //                .waitrequest
		.MASTER_READDATAVALID_AVM (traffic_gen_0_avalon_master_0_readdatavalid), //                .readdatavalid
		.MASTER_BURSTCOUNT_AVM    (traffic_gen_0_avalon_master_0_burstcount),    //                .burstcount
		.iCLOCK                   (clk_clk),                                     //      clock_sink.clk
		.iRESET                   (~rst_controller_reset_out_reset),             //      reset_sink.reset_n
		.ENABLE                   (),                                            //     conduit_end.export
		.precharge                (),                                            //                .export
		.refresh                  ()                                             //                .export
	);

	traffic_gen #(
		.SLAVE_ADDR_WIDTH  (26),
		.DATA_WIDTH        (32),
		.MASTER_ADDR_WIDTH (28),
		.BYTE_ENABLE_BITS  (4),
		.BURST_COUNT_BITS  (4),
		.BURST_LENGTH      (8),
		.NUM_OF_MASTERS    (4),
		.master_index      (1),
		.sopc_enable       (1)
	) traffic_gen_1 (
		.MASTER_ADDRES_AVM        (traffic_gen_1_avalon_master_0_address),       // avalon_master_0.address
		.MASTER_READ_AVM          (traffic_gen_1_avalon_master_0_read),          //                .read
		.MASTER_WRITE_AVM         (traffic_gen_1_avalon_master_0_write),         //                .write
		.MASTER_WRITEDATA_AVM     (traffic_gen_1_avalon_master_0_writedata),     //                .writedata
		.MASTER_BYTEENABLE_AVM    (traffic_gen_1_avalon_master_0_byteenable),    //                .byteenable
		.MASTER_READ_DATA_AVM     (traffic_gen_1_avalon_master_0_readdata),      //                .readdata
		.MASTER_WAITREQUEST_AVM   (traffic_gen_1_avalon_master_0_waitrequest),   //                .waitrequest
		.MASTER_READDATAVALID_AVM (traffic_gen_1_avalon_master_0_readdatavalid), //                .readdatavalid
		.MASTER_BURSTCOUNT_AVM    (traffic_gen_1_avalon_master_0_burstcount),    //                .burstcount
		.iCLOCK                   (clk_clk),                                     //      clock_sink.clk
		.iRESET                   (~rst_controller_reset_out_reset),             //      reset_sink.reset_n
		.ENABLE                   (),                                            //     conduit_end.export
		.precharge                (),                                            //                .export
		.refresh                  ()                                             //                .export
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (29),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (4),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (32),
		.UAV_BURSTCOUNT_W            (6),
		.USE_READ                    (1),
		.USE_WRITE                   (0),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (1),
		.USE_READDATAVALID           (1),
		.USE_WAITREQUEST             (1),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (1),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (1),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) com_nios_instruction_master_translator (
		.clk                   (clk_clk),                                                                        //                       clk.clk
		.reset                 (rst_controller_reset_out_reset),                                                 //                     reset.reset
		.uav_address           (com_nios_instruction_master_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount        (com_nios_instruction_master_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read              (com_nios_instruction_master_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write             (com_nios_instruction_master_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest       (com_nios_instruction_master_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid     (com_nios_instruction_master_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable        (com_nios_instruction_master_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata          (com_nios_instruction_master_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata         (com_nios_instruction_master_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock              (com_nios_instruction_master_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess       (com_nios_instruction_master_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address            (com_nios_instruction_master_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest        (com_nios_instruction_master_waitrequest),                                        //                          .waitrequest
		.av_burstcount         (com_nios_instruction_master_burstcount),                                         //                          .burstcount
		.av_read               (com_nios_instruction_master_read),                                               //                          .read
		.av_readdata           (com_nios_instruction_master_readdata),                                           //                          .readdata
		.av_readdatavalid      (com_nios_instruction_master_readdatavalid),                                      //                          .readdatavalid
		.av_byteenable         (4'b1111),                                                                        //               (terminated)
		.av_beginbursttransfer (1'b0),                                                                           //               (terminated)
		.av_begintransfer      (1'b0),                                                                           //               (terminated)
		.av_chipselect         (1'b0),                                                                           //               (terminated)
		.av_write              (1'b0),                                                                           //               (terminated)
		.av_writedata          (32'b00000000000000000000000000000000),                                           //               (terminated)
		.av_lock               (1'b0),                                                                           //               (terminated)
		.av_debugaccess        (1'b0),                                                                           //               (terminated)
		.uav_clken             (),                                                                               //               (terminated)
		.av_clken              (1'b1)                                                                            //               (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (29),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (4),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (32),
		.UAV_BURSTCOUNT_W            (6),
		.USE_READ                    (1),
		.USE_WRITE                   (1),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (1),
		.USE_READDATAVALID           (1),
		.USE_WAITREQUEST             (1),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (1),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) com_nios_data_master_translator (
		.clk                   (clk_clk),                                                                 //                       clk.clk
		.reset                 (rst_controller_reset_out_reset),                                          //                     reset.reset
		.uav_address           (com_nios_data_master_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount        (com_nios_data_master_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read              (com_nios_data_master_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write             (com_nios_data_master_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest       (com_nios_data_master_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid     (com_nios_data_master_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable        (com_nios_data_master_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata          (com_nios_data_master_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata         (com_nios_data_master_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock              (com_nios_data_master_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess       (com_nios_data_master_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address            (com_nios_data_master_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest        (com_nios_data_master_waitrequest),                                        //                          .waitrequest
		.av_burstcount         (com_nios_data_master_burstcount),                                         //                          .burstcount
		.av_byteenable         (com_nios_data_master_byteenable),                                         //                          .byteenable
		.av_read               (com_nios_data_master_read),                                               //                          .read
		.av_readdata           (com_nios_data_master_readdata),                                           //                          .readdata
		.av_readdatavalid      (com_nios_data_master_readdatavalid),                                      //                          .readdatavalid
		.av_write              (com_nios_data_master_write),                                              //                          .write
		.av_writedata          (com_nios_data_master_writedata),                                          //                          .writedata
		.av_debugaccess        (com_nios_data_master_debugaccess),                                        //                          .debugaccess
		.av_beginbursttransfer (1'b0),                                                                    //               (terminated)
		.av_begintransfer      (1'b0),                                                                    //               (terminated)
		.av_chipselect         (1'b0),                                                                    //               (terminated)
		.av_lock               (1'b0),                                                                    //               (terminated)
		.uav_clken             (),                                                                        //               (terminated)
		.av_clken              (1'b1)                                                                     //               (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (29),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (32),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (1),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (0),
		.USE_WAITREQUEST             (1),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) carcontrol_nios_data_master_translator (
		.clk                   (clk_clk),                                                                        //                       clk.clk
		.reset                 (rst_controller_reset_out_reset),                                                 //                     reset.reset
		.uav_address           (carcontrol_nios_data_master_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount        (carcontrol_nios_data_master_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read              (carcontrol_nios_data_master_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write             (carcontrol_nios_data_master_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest       (carcontrol_nios_data_master_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid     (carcontrol_nios_data_master_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable        (carcontrol_nios_data_master_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata          (carcontrol_nios_data_master_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata         (carcontrol_nios_data_master_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock              (carcontrol_nios_data_master_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess       (carcontrol_nios_data_master_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address            (carcontrol_nios_data_master_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest        (carcontrol_nios_data_master_waitrequest),                                        //                          .waitrequest
		.av_byteenable         (carcontrol_nios_data_master_byteenable),                                         //                          .byteenable
		.av_read               (carcontrol_nios_data_master_read),                                               //                          .read
		.av_readdata           (carcontrol_nios_data_master_readdata),                                           //                          .readdata
		.av_write              (carcontrol_nios_data_master_write),                                              //                          .write
		.av_writedata          (carcontrol_nios_data_master_writedata),                                          //                          .writedata
		.av_debugaccess        (carcontrol_nios_data_master_debugaccess),                                        //                          .debugaccess
		.av_burstcount         (1'b1),                                                                           //               (terminated)
		.av_beginbursttransfer (1'b0),                                                                           //               (terminated)
		.av_begintransfer      (1'b0),                                                                           //               (terminated)
		.av_chipselect         (1'b0),                                                                           //               (terminated)
		.av_readdatavalid      (),                                                                               //               (terminated)
		.av_lock               (1'b0),                                                                           //               (terminated)
		.uav_clken             (),                                                                               //               (terminated)
		.av_clken              (1'b1)                                                                            //               (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (29),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (32),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (0),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (1),
		.USE_WAITREQUEST             (1),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (1),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) carcontrol_nios_instruction_master_translator (
		.clk                   (clk_clk),                                                                               //                       clk.clk
		.reset                 (rst_controller_reset_out_reset),                                                        //                     reset.reset
		.uav_address           (carcontrol_nios_instruction_master_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount        (carcontrol_nios_instruction_master_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read              (carcontrol_nios_instruction_master_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write             (carcontrol_nios_instruction_master_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest       (carcontrol_nios_instruction_master_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid     (carcontrol_nios_instruction_master_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable        (carcontrol_nios_instruction_master_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata          (carcontrol_nios_instruction_master_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata         (carcontrol_nios_instruction_master_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock              (carcontrol_nios_instruction_master_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess       (carcontrol_nios_instruction_master_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address            (carcontrol_nios_instruction_master_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest        (carcontrol_nios_instruction_master_waitrequest),                                        //                          .waitrequest
		.av_read               (carcontrol_nios_instruction_master_read),                                               //                          .read
		.av_readdata           (carcontrol_nios_instruction_master_readdata),                                           //                          .readdata
		.av_readdatavalid      (carcontrol_nios_instruction_master_readdatavalid),                                      //                          .readdatavalid
		.av_burstcount         (1'b1),                                                                                  //               (terminated)
		.av_byteenable         (4'b1111),                                                                               //               (terminated)
		.av_beginbursttransfer (1'b0),                                                                                  //               (terminated)
		.av_begintransfer      (1'b0),                                                                                  //               (terminated)
		.av_chipselect         (1'b0),                                                                                  //               (terminated)
		.av_write              (1'b0),                                                                                  //               (terminated)
		.av_writedata          (32'b00000000000000000000000000000000),                                                  //               (terminated)
		.av_lock               (1'b0),                                                                                  //               (terminated)
		.av_debugaccess        (1'b0),                                                                                  //               (terminated)
		.uav_clken             (),                                                                                      //               (terminated)
		.av_clken              (1'b1)                                                                                   //               (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (32),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (32),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (0),
		.USE_WRITE                   (1),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (0),
		.USE_WAITREQUEST             (1),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) ethernet_subsystem_sgdma_rx_m_write_translator (
		.clk                   (clk_clk),                                                                                //                       clk.clk
		.reset                 (rst_controller_002_reset_out_reset),                                                     //                     reset.reset
		.uav_address           (ethernet_subsystem_sgdma_rx_m_write_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount        (ethernet_subsystem_sgdma_rx_m_write_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read              (ethernet_subsystem_sgdma_rx_m_write_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write             (ethernet_subsystem_sgdma_rx_m_write_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest       (ethernet_subsystem_sgdma_rx_m_write_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid     (ethernet_subsystem_sgdma_rx_m_write_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable        (ethernet_subsystem_sgdma_rx_m_write_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata          (ethernet_subsystem_sgdma_rx_m_write_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata         (ethernet_subsystem_sgdma_rx_m_write_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock              (ethernet_subsystem_sgdma_rx_m_write_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess       (ethernet_subsystem_sgdma_rx_m_write_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address            (ethernet_subsystem_sgdma_rx_m_write_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest        (ethernet_subsystem_sgdma_rx_m_write_waitrequest),                                        //                          .waitrequest
		.av_byteenable         (ethernet_subsystem_sgdma_rx_m_write_byteenable),                                         //                          .byteenable
		.av_write              (ethernet_subsystem_sgdma_rx_m_write_write),                                              //                          .write
		.av_writedata          (ethernet_subsystem_sgdma_rx_m_write_writedata),                                          //                          .writedata
		.av_burstcount         (1'b1),                                                                                   //               (terminated)
		.av_beginbursttransfer (1'b0),                                                                                   //               (terminated)
		.av_begintransfer      (1'b0),                                                                                   //               (terminated)
		.av_chipselect         (1'b0),                                                                                   //               (terminated)
		.av_read               (1'b0),                                                                                   //               (terminated)
		.av_readdata           (),                                                                                       //               (terminated)
		.av_readdatavalid      (),                                                                                       //               (terminated)
		.av_lock               (1'b0),                                                                                   //               (terminated)
		.av_debugaccess        (1'b0),                                                                                   //               (terminated)
		.uav_clken             (),                                                                                       //               (terminated)
		.av_clken              (1'b1)                                                                                    //               (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (32),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (32),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (0),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (1),
		.USE_WAITREQUEST             (1),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) ethernet_subsystem_sgdma_tx_m_read_translator (
		.clk                   (clk_clk),                                                                               //                       clk.clk
		.reset                 (rst_controller_002_reset_out_reset),                                                    //                     reset.reset
		.uav_address           (ethernet_subsystem_sgdma_tx_m_read_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount        (ethernet_subsystem_sgdma_tx_m_read_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read              (ethernet_subsystem_sgdma_tx_m_read_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write             (ethernet_subsystem_sgdma_tx_m_read_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest       (ethernet_subsystem_sgdma_tx_m_read_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid     (ethernet_subsystem_sgdma_tx_m_read_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable        (ethernet_subsystem_sgdma_tx_m_read_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata          (ethernet_subsystem_sgdma_tx_m_read_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata         (ethernet_subsystem_sgdma_tx_m_read_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock              (ethernet_subsystem_sgdma_tx_m_read_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess       (ethernet_subsystem_sgdma_tx_m_read_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address            (ethernet_subsystem_sgdma_tx_m_read_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest        (ethernet_subsystem_sgdma_tx_m_read_waitrequest),                                        //                          .waitrequest
		.av_read               (ethernet_subsystem_sgdma_tx_m_read_read),                                               //                          .read
		.av_readdata           (ethernet_subsystem_sgdma_tx_m_read_readdata),                                           //                          .readdata
		.av_readdatavalid      (ethernet_subsystem_sgdma_tx_m_read_readdatavalid),                                      //                          .readdatavalid
		.av_burstcount         (1'b1),                                                                                  //               (terminated)
		.av_byteenable         (4'b1111),                                                                               //               (terminated)
		.av_beginbursttransfer (1'b0),                                                                                  //               (terminated)
		.av_begintransfer      (1'b0),                                                                                  //               (terminated)
		.av_chipselect         (1'b0),                                                                                  //               (terminated)
		.av_write              (1'b0),                                                                                  //               (terminated)
		.av_writedata          (32'b00000000000000000000000000000000),                                                  //               (terminated)
		.av_lock               (1'b0),                                                                                  //               (terminated)
		.av_debugaccess        (1'b0),                                                                                  //               (terminated)
		.uav_clken             (),                                                                                      //               (terminated)
		.av_clken              (1'b1)                                                                                   //               (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (9),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) com_nios_jtag_debug_module_translator (
		.clk                   (clk_clk),                                                                               //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                                        //                    reset.reset
		.uav_address           (com_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (com_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (com_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (com_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (com_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (com_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (com_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (com_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (com_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (com_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (com_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (com_nios_jtag_debug_module_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (com_nios_jtag_debug_module_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (com_nios_jtag_debug_module_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (com_nios_jtag_debug_module_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_begintransfer      (com_nios_jtag_debug_module_translator_avalon_anti_slave_0_begintransfer),               //                         .begintransfer
		.av_byteenable         (com_nios_jtag_debug_module_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_chipselect         (com_nios_jtag_debug_module_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_debugaccess        (com_nios_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess),                 //                         .debugaccess
		.av_read               (),                                                                                      //              (terminated)
		.av_beginbursttransfer (),                                                                                      //              (terminated)
		.av_burstcount         (),                                                                                      //              (terminated)
		.av_readdatavalid      (1'b0),                                                                                  //              (terminated)
		.av_waitrequest        (1'b0),                                                                                  //              (terminated)
		.av_writebyteenable    (),                                                                                      //              (terminated)
		.av_lock               (),                                                                                      //              (terminated)
		.av_clken              (),                                                                                      //              (terminated)
		.uav_clken             (1'b0),                                                                                  //              (terminated)
		.av_outputenable       ()                                                                                       //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (24),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (1),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) com_memory_s1_translator (
		.clk                   (clk_clk),                                                                  //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                           //                    reset.reset
		.uav_address           (com_memory_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (com_memory_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (com_memory_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (com_memory_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (com_memory_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (com_memory_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (com_memory_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (com_memory_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (com_memory_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (com_memory_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (com_memory_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (com_memory_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (com_memory_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (com_memory_s1_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (com_memory_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (com_memory_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable         (com_memory_s1_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_readdatavalid      (com_memory_s1_translator_avalon_anti_slave_0_readdatavalid),               //                         .readdatavalid
		.av_waitrequest        (com_memory_s1_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_chipselect         (com_memory_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer      (),                                                                         //              (terminated)
		.av_beginbursttransfer (),                                                                         //              (terminated)
		.av_burstcount         (),                                                                         //              (terminated)
		.av_writebyteenable    (),                                                                         //              (terminated)
		.av_lock               (),                                                                         //              (terminated)
		.av_clken              (),                                                                         //              (terminated)
		.uav_clken             (1'b0),                                                                     //              (terminated)
		.av_debugaccess        (),                                                                         //              (terminated)
		.av_outputenable       ()                                                                          //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) jtaguart_0_avalon_jtag_slave_translator (
		.clk                   (clk_clk),                                                                                 //                      clk.clk
		.reset                 (rst_controller_001_reset_out_reset),                                                      //                    reset.reset
		.uav_address           (jtaguart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (jtaguart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (jtaguart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (jtaguart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (jtaguart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (jtaguart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (jtaguart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (jtaguart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (jtaguart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (jtaguart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (jtaguart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (jtaguart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (jtaguart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (jtaguart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (jtaguart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (jtaguart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_waitrequest        (jtaguart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_chipselect         (jtaguart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer      (),                                                                                        //              (terminated)
		.av_beginbursttransfer (),                                                                                        //              (terminated)
		.av_burstcount         (),                                                                                        //              (terminated)
		.av_byteenable         (),                                                                                        //              (terminated)
		.av_readdatavalid      (1'b0),                                                                                    //              (terminated)
		.av_writebyteenable    (),                                                                                        //              (terminated)
		.av_lock               (),                                                                                        //              (terminated)
		.av_clken              (),                                                                                        //              (terminated)
		.uav_clken             (1'b0),                                                                                    //              (terminated)
		.av_debugaccess        (),                                                                                        //              (terminated)
		.av_outputenable       ()                                                                                         //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) shared_memory_mutex_s1_translator (
		.clk                   (clk_clk),                                                                           //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                                    //                    reset.reset
		.uav_address           (shared_memory_mutex_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (shared_memory_mutex_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (shared_memory_mutex_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (shared_memory_mutex_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (shared_memory_mutex_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (shared_memory_mutex_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (shared_memory_mutex_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (shared_memory_mutex_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (shared_memory_mutex_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (shared_memory_mutex_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (shared_memory_mutex_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (shared_memory_mutex_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (shared_memory_mutex_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (shared_memory_mutex_s1_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (shared_memory_mutex_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (shared_memory_mutex_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect         (shared_memory_mutex_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer      (),                                                                                  //              (terminated)
		.av_beginbursttransfer (),                                                                                  //              (terminated)
		.av_burstcount         (),                                                                                  //              (terminated)
		.av_byteenable         (),                                                                                  //              (terminated)
		.av_readdatavalid      (1'b0),                                                                              //              (terminated)
		.av_waitrequest        (1'b0),                                                                              //              (terminated)
		.av_writebyteenable    (),                                                                                  //              (terminated)
		.av_lock               (),                                                                                  //              (terminated)
		.av_clken              (),                                                                                  //              (terminated)
		.uav_clken             (1'b0),                                                                              //              (terminated)
		.av_debugaccess        (),                                                                                  //              (terminated)
		.av_outputenable       ()                                                                                   //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (3),
		.AV_DATA_W                      (16),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) com_timer_s1_translator (
		.clk                   (clk_clk),                                                                 //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                          //                    reset.reset
		.uav_address           (com_timer_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (com_timer_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (com_timer_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (com_timer_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (com_timer_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (com_timer_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (com_timer_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (com_timer_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (com_timer_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (com_timer_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (com_timer_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (com_timer_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (com_timer_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (com_timer_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (com_timer_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect         (com_timer_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read               (),                                                                        //              (terminated)
		.av_begintransfer      (),                                                                        //              (terminated)
		.av_beginbursttransfer (),                                                                        //              (terminated)
		.av_burstcount         (),                                                                        //              (terminated)
		.av_byteenable         (),                                                                        //              (terminated)
		.av_readdatavalid      (1'b0),                                                                    //              (terminated)
		.av_waitrequest        (1'b0),                                                                    //              (terminated)
		.av_writebyteenable    (),                                                                        //              (terminated)
		.av_lock               (),                                                                        //              (terminated)
		.av_clken              (),                                                                        //              (terminated)
		.uav_clken             (1'b0),                                                                    //              (terminated)
		.av_debugaccess        (),                                                                        //              (terminated)
		.av_outputenable       ()                                                                         //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (11),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (1),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (1),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) ethernet_subsystem_ethernet_bridge_s0_translator (
		.clk                   (clk_clk),                                                                                          //                      clk.clk
		.reset                 (rst_controller_002_reset_out_reset),                                                               //                    reset.reset
		.uav_address           (ethernet_subsystem_ethernet_bridge_s0_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (ethernet_subsystem_ethernet_bridge_s0_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (ethernet_subsystem_ethernet_bridge_s0_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (ethernet_subsystem_ethernet_bridge_s0_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (ethernet_subsystem_ethernet_bridge_s0_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (ethernet_subsystem_ethernet_bridge_s0_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (ethernet_subsystem_ethernet_bridge_s0_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (ethernet_subsystem_ethernet_bridge_s0_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (ethernet_subsystem_ethernet_bridge_s0_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (ethernet_subsystem_ethernet_bridge_s0_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (ethernet_subsystem_ethernet_bridge_s0_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (ethernet_subsystem_ethernet_bridge_s0_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (ethernet_subsystem_ethernet_bridge_s0_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (ethernet_subsystem_ethernet_bridge_s0_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (ethernet_subsystem_ethernet_bridge_s0_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (ethernet_subsystem_ethernet_bridge_s0_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_burstcount         (ethernet_subsystem_ethernet_bridge_s0_translator_avalon_anti_slave_0_burstcount),                  //                         .burstcount
		.av_byteenable         (ethernet_subsystem_ethernet_bridge_s0_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_readdatavalid      (ethernet_subsystem_ethernet_bridge_s0_translator_avalon_anti_slave_0_readdatavalid),               //                         .readdatavalid
		.av_waitrequest        (ethernet_subsystem_ethernet_bridge_s0_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_debugaccess        (ethernet_subsystem_ethernet_bridge_s0_translator_avalon_anti_slave_0_debugaccess),                 //                         .debugaccess
		.av_begintransfer      (),                                                                                                 //              (terminated)
		.av_beginbursttransfer (),                                                                                                 //              (terminated)
		.av_writebyteenable    (),                                                                                                 //              (terminated)
		.av_lock               (),                                                                                                 //              (terminated)
		.av_chipselect         (),                                                                                                 //              (terminated)
		.av_clken              (),                                                                                                 //              (terminated)
		.uav_clken             (1'b0),                                                                                             //              (terminated)
		.av_outputenable       ()                                                                                                  //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (11),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (1),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) ethernet_subsystem_descriptor_memory_s2_translator (
		.clk                   (clk_clk),                                                                                            //                      clk.clk
		.reset                 (rst_controller_002_reset_out_reset),                                                                 //                    reset.reset
		.uav_address           (ethernet_subsystem_descriptor_memory_s2_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (ethernet_subsystem_descriptor_memory_s2_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (ethernet_subsystem_descriptor_memory_s2_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (ethernet_subsystem_descriptor_memory_s2_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (ethernet_subsystem_descriptor_memory_s2_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (ethernet_subsystem_descriptor_memory_s2_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (ethernet_subsystem_descriptor_memory_s2_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (ethernet_subsystem_descriptor_memory_s2_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (ethernet_subsystem_descriptor_memory_s2_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (ethernet_subsystem_descriptor_memory_s2_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (ethernet_subsystem_descriptor_memory_s2_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (ethernet_subsystem_descriptor_memory_s2_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (ethernet_subsystem_descriptor_memory_s2_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (ethernet_subsystem_descriptor_memory_s2_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (ethernet_subsystem_descriptor_memory_s2_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable         (ethernet_subsystem_descriptor_memory_s2_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_chipselect         (ethernet_subsystem_descriptor_memory_s2_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_clken              (ethernet_subsystem_descriptor_memory_s2_translator_avalon_anti_slave_0_clken),                       //                         .clken
		.av_read               (),                                                                                                   //              (terminated)
		.av_begintransfer      (),                                                                                                   //              (terminated)
		.av_beginbursttransfer (),                                                                                                   //              (terminated)
		.av_burstcount         (),                                                                                                   //              (terminated)
		.av_readdatavalid      (1'b0),                                                                                               //              (terminated)
		.av_waitrequest        (1'b0),                                                                                               //              (terminated)
		.av_writebyteenable    (),                                                                                                   //              (terminated)
		.av_lock               (),                                                                                                   //              (terminated)
		.uav_clken             (1'b0),                                                                                               //              (terminated)
		.av_debugaccess        (),                                                                                                   //              (terminated)
		.av_outputenable       ()                                                                                                    //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (26),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (1),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) prio_arbiter_0_s0_translator (
		.clk                   (clk_clk),                                                                      //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                               //                    reset.reset
		.uav_address           (prio_arbiter_0_s0_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (prio_arbiter_0_s0_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (prio_arbiter_0_s0_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (prio_arbiter_0_s0_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (prio_arbiter_0_s0_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (prio_arbiter_0_s0_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (prio_arbiter_0_s0_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (prio_arbiter_0_s0_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (prio_arbiter_0_s0_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (prio_arbiter_0_s0_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (prio_arbiter_0_s0_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (prio_arbiter_0_s0_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (prio_arbiter_0_s0_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (prio_arbiter_0_s0_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (prio_arbiter_0_s0_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (prio_arbiter_0_s0_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable         (prio_arbiter_0_s0_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_readdatavalid      (prio_arbiter_0_s0_translator_avalon_anti_slave_0_readdatavalid),               //                         .readdatavalid
		.av_waitrequest        (prio_arbiter_0_s0_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_chipselect         (prio_arbiter_0_s0_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer      (),                                                                             //              (terminated)
		.av_beginbursttransfer (),                                                                             //              (terminated)
		.av_burstcount         (),                                                                             //              (terminated)
		.av_writebyteenable    (),                                                                             //              (terminated)
		.av_lock               (),                                                                             //              (terminated)
		.av_clken              (),                                                                             //              (terminated)
		.uav_clken             (1'b0),                                                                         //              (terminated)
		.av_debugaccess        (),                                                                             //              (terminated)
		.av_outputenable       ()                                                                              //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (9),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) carcontrol_nios_jtag_debug_module_translator (
		.clk                   (clk_clk),                                                                                      //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                                               //                    reset.reset
		.uav_address           (carcontrol_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (carcontrol_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (carcontrol_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (carcontrol_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (carcontrol_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (carcontrol_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (carcontrol_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (carcontrol_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (carcontrol_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (carcontrol_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (carcontrol_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (carcontrol_nios_jtag_debug_module_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (carcontrol_nios_jtag_debug_module_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (carcontrol_nios_jtag_debug_module_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (carcontrol_nios_jtag_debug_module_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_begintransfer      (carcontrol_nios_jtag_debug_module_translator_avalon_anti_slave_0_begintransfer),               //                         .begintransfer
		.av_byteenable         (carcontrol_nios_jtag_debug_module_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_chipselect         (carcontrol_nios_jtag_debug_module_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_debugaccess        (carcontrol_nios_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess),                 //                         .debugaccess
		.av_read               (),                                                                                             //              (terminated)
		.av_beginbursttransfer (),                                                                                             //              (terminated)
		.av_burstcount         (),                                                                                             //              (terminated)
		.av_readdatavalid      (1'b0),                                                                                         //              (terminated)
		.av_waitrequest        (1'b0),                                                                                         //              (terminated)
		.av_writebyteenable    (),                                                                                             //              (terminated)
		.av_lock               (),                                                                                             //              (terminated)
		.av_clken              (),                                                                                             //              (terminated)
		.uav_clken             (1'b0),                                                                                         //              (terminated)
		.av_outputenable       ()                                                                                              //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (16),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (1),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) onchip_memory2_0_s1_translator (
		.clk                   (clk_clk),                                                                        //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                                 //                    reset.reset
		.uav_address           (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (onchip_memory2_0_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (onchip_memory2_0_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (onchip_memory2_0_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (onchip_memory2_0_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable         (onchip_memory2_0_s1_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_chipselect         (onchip_memory2_0_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_clken              (onchip_memory2_0_s1_translator_avalon_anti_slave_0_clken),                       //                         .clken
		.av_read               (),                                                                               //              (terminated)
		.av_begintransfer      (),                                                                               //              (terminated)
		.av_beginbursttransfer (),                                                                               //              (terminated)
		.av_burstcount         (),                                                                               //              (terminated)
		.av_readdatavalid      (1'b0),                                                                           //              (terminated)
		.av_waitrequest        (1'b0),                                                                           //              (terminated)
		.av_writebyteenable    (),                                                                               //              (terminated)
		.av_lock               (),                                                                               //              (terminated)
		.uav_clken             (1'b0),                                                                           //              (terminated)
		.av_debugaccess        (),                                                                               //              (terminated)
		.av_outputenable       ()                                                                                //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) jtaguart_1_avalon_jtag_slave_translator (
		.clk                   (clk_clk),                                                                                 //                      clk.clk
		.reset                 (rst_controller_002_reset_out_reset),                                                      //                    reset.reset
		.uav_address           (jtaguart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (jtaguart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (jtaguart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (jtaguart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (jtaguart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (jtaguart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (jtaguart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (jtaguart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (jtaguart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (jtaguart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (jtaguart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (jtaguart_1_avalon_jtag_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (jtaguart_1_avalon_jtag_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (jtaguart_1_avalon_jtag_slave_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (jtaguart_1_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (jtaguart_1_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_waitrequest        (jtaguart_1_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_chipselect         (jtaguart_1_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer      (),                                                                                        //              (terminated)
		.av_beginbursttransfer (),                                                                                        //              (terminated)
		.av_burstcount         (),                                                                                        //              (terminated)
		.av_byteenable         (),                                                                                        //              (terminated)
		.av_readdatavalid      (1'b0),                                                                                    //              (terminated)
		.av_writebyteenable    (),                                                                                        //              (terminated)
		.av_lock               (),                                                                                        //              (terminated)
		.av_clken              (),                                                                                        //              (terminated)
		.uav_clken             (1'b0),                                                                                    //              (terminated)
		.av_debugaccess        (),                                                                                        //              (terminated)
		.av_outputenable       ()                                                                                         //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (26),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (1),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) prio_arbiter_0_s1_translator (
		.clk                   (clk_clk),                                                                      //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                               //                    reset.reset
		.uav_address           (prio_arbiter_0_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (prio_arbiter_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (prio_arbiter_0_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (prio_arbiter_0_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (prio_arbiter_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (prio_arbiter_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (prio_arbiter_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (prio_arbiter_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (prio_arbiter_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (prio_arbiter_0_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (prio_arbiter_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (prio_arbiter_0_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (prio_arbiter_0_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (prio_arbiter_0_s1_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (prio_arbiter_0_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (prio_arbiter_0_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable         (prio_arbiter_0_s1_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_readdatavalid      (prio_arbiter_0_s1_translator_avalon_anti_slave_0_readdatavalid),               //                         .readdatavalid
		.av_waitrequest        (prio_arbiter_0_s1_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_chipselect         (prio_arbiter_0_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer      (),                                                                             //              (terminated)
		.av_beginbursttransfer (),                                                                             //              (terminated)
		.av_burstcount         (),                                                                             //              (terminated)
		.av_writebyteenable    (),                                                                             //              (terminated)
		.av_lock               (),                                                                             //              (terminated)
		.av_clken              (),                                                                             //              (terminated)
		.uav_clken             (1'b0),                                                                         //              (terminated)
		.av_debugaccess        (),                                                                             //              (terminated)
		.av_outputenable       ()                                                                              //              (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (28),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (28),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (1),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (1),
		.USE_WAITREQUEST             (1),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) prio_arbiter_0_m1_translator (
		.clk                   (clk_clk),                                                              //                       clk.clk
		.reset                 (rst_controller_reset_out_reset),                                       //                     reset.reset
		.uav_address           (prio_arbiter_0_m1_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount        (prio_arbiter_0_m1_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read              (prio_arbiter_0_m1_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write             (prio_arbiter_0_m1_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest       (prio_arbiter_0_m1_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid     (prio_arbiter_0_m1_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable        (prio_arbiter_0_m1_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata          (prio_arbiter_0_m1_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata         (prio_arbiter_0_m1_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock              (prio_arbiter_0_m1_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess       (prio_arbiter_0_m1_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address            (prio_arbiter_0_m1_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest        (prio_arbiter_0_m1_waitrequest),                                        //                          .waitrequest
		.av_byteenable         (prio_arbiter_0_m1_byteenable),                                         //                          .byteenable
		.av_read               (prio_arbiter_0_m1_read),                                               //                          .read
		.av_readdata           (prio_arbiter_0_m1_readdata),                                           //                          .readdata
		.av_readdatavalid      (prio_arbiter_0_m1_readdatavalid),                                      //                          .readdatavalid
		.av_write              (prio_arbiter_0_m1_write),                                              //                          .write
		.av_writedata          (prio_arbiter_0_m1_writedata),                                          //                          .writedata
		.av_burstcount         (1'b1),                                                                 //               (terminated)
		.av_beginbursttransfer (1'b0),                                                                 //               (terminated)
		.av_begintransfer      (1'b0),                                                                 //               (terminated)
		.av_chipselect         (1'b0),                                                                 //               (terminated)
		.av_lock               (1'b0),                                                                 //               (terminated)
		.av_debugaccess        (1'b0),                                                                 //               (terminated)
		.uav_clken             (),                                                                     //               (terminated)
		.av_clken              (1'b1)                                                                  //               (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (10),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (28),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (1),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) shared_memory_s1_translator (
		.clk                   (clk_clk),                                                              //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                       //                    reset.reset
		.uav_address           (prio_arbiter_0_m1_translator_avalon_universal_master_0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (prio_arbiter_0_m1_translator_avalon_universal_master_0_burstcount),    //                         .burstcount
		.uav_read              (prio_arbiter_0_m1_translator_avalon_universal_master_0_read),          //                         .read
		.uav_write             (prio_arbiter_0_m1_translator_avalon_universal_master_0_write),         //                         .write
		.uav_waitrequest       (prio_arbiter_0_m1_translator_avalon_universal_master_0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (prio_arbiter_0_m1_translator_avalon_universal_master_0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (prio_arbiter_0_m1_translator_avalon_universal_master_0_byteenable),    //                         .byteenable
		.uav_readdata          (prio_arbiter_0_m1_translator_avalon_universal_master_0_readdata),      //                         .readdata
		.uav_writedata         (prio_arbiter_0_m1_translator_avalon_universal_master_0_writedata),     //                         .writedata
		.uav_lock              (prio_arbiter_0_m1_translator_avalon_universal_master_0_lock),          //                         .lock
		.uav_debugaccess       (prio_arbiter_0_m1_translator_avalon_universal_master_0_debugaccess),   //                         .debugaccess
		.av_address            (shared_memory_s1_translator_avalon_anti_slave_0_address),              //      avalon_anti_slave_0.address
		.av_write              (shared_memory_s1_translator_avalon_anti_slave_0_write),                //                         .write
		.av_readdata           (shared_memory_s1_translator_avalon_anti_slave_0_readdata),             //                         .readdata
		.av_writedata          (shared_memory_s1_translator_avalon_anti_slave_0_writedata),            //                         .writedata
		.av_byteenable         (shared_memory_s1_translator_avalon_anti_slave_0_byteenable),           //                         .byteenable
		.av_chipselect         (shared_memory_s1_translator_avalon_anti_slave_0_chipselect),           //                         .chipselect
		.av_clken              (shared_memory_s1_translator_avalon_anti_slave_0_clken),                //                         .clken
		.av_read               (),                                                                     //              (terminated)
		.av_begintransfer      (),                                                                     //              (terminated)
		.av_beginbursttransfer (),                                                                     //              (terminated)
		.av_burstcount         (),                                                                     //              (terminated)
		.av_readdatavalid      (1'b0),                                                                 //              (terminated)
		.av_waitrequest        (1'b0),                                                                 //              (terminated)
		.av_writebyteenable    (),                                                                     //              (terminated)
		.av_lock               (),                                                                     //              (terminated)
		.uav_clken             (1'b0),                                                                 //              (terminated)
		.av_debugaccess        (),                                                                     //              (terminated)
		.av_outputenable       ()                                                                      //              (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (28),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (4),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (28),
		.UAV_BURSTCOUNT_W            (6),
		.USE_READ                    (1),
		.USE_WRITE                   (1),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (1),
		.USE_READDATAVALID           (1),
		.USE_WAITREQUEST             (1),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (1),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) traffic_gen_0_avalon_master_0_translator (
		.clk                   (clk_clk),                                                                          //                       clk.clk
		.reset                 (rst_controller_reset_out_reset),                                                   //                     reset.reset
		.uav_address           (traffic_gen_0_avalon_master_0_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount        (traffic_gen_0_avalon_master_0_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read              (traffic_gen_0_avalon_master_0_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write             (traffic_gen_0_avalon_master_0_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest       (traffic_gen_0_avalon_master_0_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid     (traffic_gen_0_avalon_master_0_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable        (traffic_gen_0_avalon_master_0_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata          (traffic_gen_0_avalon_master_0_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata         (traffic_gen_0_avalon_master_0_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock              (traffic_gen_0_avalon_master_0_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess       (traffic_gen_0_avalon_master_0_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address            (traffic_gen_0_avalon_master_0_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest        (traffic_gen_0_avalon_master_0_waitrequest),                                        //                          .waitrequest
		.av_burstcount         (traffic_gen_0_avalon_master_0_burstcount),                                         //                          .burstcount
		.av_byteenable         (traffic_gen_0_avalon_master_0_byteenable),                                         //                          .byteenable
		.av_read               (traffic_gen_0_avalon_master_0_read),                                               //                          .read
		.av_readdata           (traffic_gen_0_avalon_master_0_readdata),                                           //                          .readdata
		.av_readdatavalid      (traffic_gen_0_avalon_master_0_readdatavalid),                                      //                          .readdatavalid
		.av_write              (traffic_gen_0_avalon_master_0_write),                                              //                          .write
		.av_writedata          (traffic_gen_0_avalon_master_0_writedata),                                          //                          .writedata
		.av_beginbursttransfer (1'b0),                                                                             //               (terminated)
		.av_begintransfer      (1'b0),                                                                             //               (terminated)
		.av_chipselect         (1'b0),                                                                             //               (terminated)
		.av_lock               (1'b0),                                                                             //               (terminated)
		.av_debugaccess        (1'b0),                                                                             //               (terminated)
		.uav_clken             (),                                                                                 //               (terminated)
		.av_clken              (1'b1)                                                                              //               (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (26),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (28),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (1),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) prio_arbiter_0_s2_translator (
		.clk                   (clk_clk),                                                                      //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                               //                    reset.reset
		.uav_address           (prio_arbiter_0_s2_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (prio_arbiter_0_s2_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (prio_arbiter_0_s2_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (prio_arbiter_0_s2_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (prio_arbiter_0_s2_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (prio_arbiter_0_s2_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (prio_arbiter_0_s2_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (prio_arbiter_0_s2_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (prio_arbiter_0_s2_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (prio_arbiter_0_s2_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (prio_arbiter_0_s2_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (prio_arbiter_0_s2_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (prio_arbiter_0_s2_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (prio_arbiter_0_s2_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (prio_arbiter_0_s2_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (prio_arbiter_0_s2_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable         (prio_arbiter_0_s2_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_readdatavalid      (prio_arbiter_0_s2_translator_avalon_anti_slave_0_readdatavalid),               //                         .readdatavalid
		.av_waitrequest        (prio_arbiter_0_s2_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_chipselect         (prio_arbiter_0_s2_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer      (),                                                                             //              (terminated)
		.av_beginbursttransfer (),                                                                             //              (terminated)
		.av_burstcount         (),                                                                             //              (terminated)
		.av_writebyteenable    (),                                                                             //              (terminated)
		.av_lock               (),                                                                             //              (terminated)
		.av_clken              (),                                                                             //              (terminated)
		.uav_clken             (1'b0),                                                                         //              (terminated)
		.av_debugaccess        (),                                                                             //              (terminated)
		.av_outputenable       ()                                                                              //              (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (28),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (4),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (28),
		.UAV_BURSTCOUNT_W            (6),
		.USE_READ                    (1),
		.USE_WRITE                   (1),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (1),
		.USE_READDATAVALID           (1),
		.USE_WAITREQUEST             (1),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (1),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) traffic_gen_1_avalon_master_0_translator (
		.clk                   (clk_clk),                                                                          //                       clk.clk
		.reset                 (rst_controller_reset_out_reset),                                                   //                     reset.reset
		.uav_address           (traffic_gen_1_avalon_master_0_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount        (traffic_gen_1_avalon_master_0_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read              (traffic_gen_1_avalon_master_0_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write             (traffic_gen_1_avalon_master_0_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest       (traffic_gen_1_avalon_master_0_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid     (traffic_gen_1_avalon_master_0_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable        (traffic_gen_1_avalon_master_0_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata          (traffic_gen_1_avalon_master_0_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata         (traffic_gen_1_avalon_master_0_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock              (traffic_gen_1_avalon_master_0_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess       (traffic_gen_1_avalon_master_0_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address            (traffic_gen_1_avalon_master_0_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest        (traffic_gen_1_avalon_master_0_waitrequest),                                        //                          .waitrequest
		.av_burstcount         (traffic_gen_1_avalon_master_0_burstcount),                                         //                          .burstcount
		.av_byteenable         (traffic_gen_1_avalon_master_0_byteenable),                                         //                          .byteenable
		.av_read               (traffic_gen_1_avalon_master_0_read),                                               //                          .read
		.av_readdata           (traffic_gen_1_avalon_master_0_readdata),                                           //                          .readdata
		.av_readdatavalid      (traffic_gen_1_avalon_master_0_readdatavalid),                                      //                          .readdatavalid
		.av_write              (traffic_gen_1_avalon_master_0_write),                                              //                          .write
		.av_writedata          (traffic_gen_1_avalon_master_0_writedata),                                          //                          .writedata
		.av_beginbursttransfer (1'b0),                                                                             //               (terminated)
		.av_begintransfer      (1'b0),                                                                             //               (terminated)
		.av_chipselect         (1'b0),                                                                             //               (terminated)
		.av_lock               (1'b0),                                                                             //               (terminated)
		.av_debugaccess        (1'b0),                                                                             //               (terminated)
		.uav_clken             (),                                                                                 //               (terminated)
		.av_clken              (1'b1)                                                                              //               (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (26),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (28),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (1),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) prio_arbiter_0_s3_translator (
		.clk                   (clk_clk),                                                                      //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                               //                    reset.reset
		.uav_address           (prio_arbiter_0_s3_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (prio_arbiter_0_s3_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (prio_arbiter_0_s3_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (prio_arbiter_0_s3_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (prio_arbiter_0_s3_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (prio_arbiter_0_s3_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (prio_arbiter_0_s3_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (prio_arbiter_0_s3_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (prio_arbiter_0_s3_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (prio_arbiter_0_s3_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (prio_arbiter_0_s3_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (prio_arbiter_0_s3_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (prio_arbiter_0_s3_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (prio_arbiter_0_s3_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (prio_arbiter_0_s3_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (prio_arbiter_0_s3_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable         (prio_arbiter_0_s3_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_readdatavalid      (prio_arbiter_0_s3_translator_avalon_anti_slave_0_readdatavalid),               //                         .readdatavalid
		.av_waitrequest        (prio_arbiter_0_s3_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_chipselect         (prio_arbiter_0_s3_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer      (),                                                                             //              (terminated)
		.av_beginbursttransfer (),                                                                             //              (terminated)
		.av_burstcount         (),                                                                             //              (terminated)
		.av_writebyteenable    (),                                                                             //              (terminated)
		.av_lock               (),                                                                             //              (terminated)
		.av_clken              (),                                                                             //              (terminated)
		.uav_clken             (1'b0),                                                                         //              (terminated)
		.av_debugaccess        (),                                                                             //              (terminated)
		.av_outputenable       ()                                                                              //              (terminated)
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (106),
		.PKT_PROTECTION_L          (104),
		.PKT_BEGIN_BURST           (93),
		.PKT_BURSTWRAP_H           (85),
		.PKT_BURSTWRAP_L           (80),
		.PKT_BURST_SIZE_H          (88),
		.PKT_BURST_SIZE_L          (86),
		.PKT_BURST_TYPE_H          (90),
		.PKT_BURST_TYPE_L          (89),
		.PKT_BYTE_CNT_H            (79),
		.PKT_BYTE_CNT_L            (74),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_TRANS_EXCLUSIVE       (73),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (98),
		.PKT_SRC_ID_L              (95),
		.PKT_DEST_ID_H             (102),
		.PKT_DEST_ID_L             (99),
		.PKT_THREAD_ID_H           (103),
		.PKT_THREAD_ID_L           (103),
		.PKT_CACHE_H               (110),
		.PKT_CACHE_L               (107),
		.PKT_DATA_SIDEBAND_H       (92),
		.PKT_DATA_SIDEBAND_L       (92),
		.PKT_QOS_H                 (94),
		.PKT_QOS_L                 (94),
		.PKT_ADDR_SIDEBAND_H       (91),
		.PKT_ADDR_SIDEBAND_L       (91),
		.ST_DATA_W                 (113),
		.ST_CHANNEL_W              (12),
		.AV_BURSTCOUNT_W           (6),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (0),
		.BURSTWRAP_VALUE           (31),
		.CACHE_VALUE               (4'b0000)
	) com_nios_instruction_master_translator_avalon_universal_master_0_agent (
		.clk              (clk_clk),                                                                                 //       clk.clk
		.reset            (rst_controller_reset_out_reset),                                                          // clk_reset.reset
		.av_address       (com_nios_instruction_master_translator_avalon_universal_master_0_address),                //        av.address
		.av_write         (com_nios_instruction_master_translator_avalon_universal_master_0_write),                  //          .write
		.av_read          (com_nios_instruction_master_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata     (com_nios_instruction_master_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata      (com_nios_instruction_master_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest   (com_nios_instruction_master_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid (com_nios_instruction_master_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable    (com_nios_instruction_master_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount    (com_nios_instruction_master_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess   (com_nios_instruction_master_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock          (com_nios_instruction_master_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid         (com_nios_instruction_master_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data          (com_nios_instruction_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket (com_nios_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket   (com_nios_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready         (com_nios_instruction_master_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid         (limiter_rsp_src_valid),                                                                   //        rp.valid
		.rp_data          (limiter_rsp_src_data),                                                                    //          .data
		.rp_channel       (limiter_rsp_src_channel),                                                                 //          .channel
		.rp_startofpacket (limiter_rsp_src_startofpacket),                                                           //          .startofpacket
		.rp_endofpacket   (limiter_rsp_src_endofpacket),                                                             //          .endofpacket
		.rp_ready         (limiter_rsp_src_ready)                                                                    //          .ready
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (106),
		.PKT_PROTECTION_L          (104),
		.PKT_BEGIN_BURST           (93),
		.PKT_BURSTWRAP_H           (85),
		.PKT_BURSTWRAP_L           (80),
		.PKT_BURST_SIZE_H          (88),
		.PKT_BURST_SIZE_L          (86),
		.PKT_BURST_TYPE_H          (90),
		.PKT_BURST_TYPE_L          (89),
		.PKT_BYTE_CNT_H            (79),
		.PKT_BYTE_CNT_L            (74),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_TRANS_EXCLUSIVE       (73),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (98),
		.PKT_SRC_ID_L              (95),
		.PKT_DEST_ID_H             (102),
		.PKT_DEST_ID_L             (99),
		.PKT_THREAD_ID_H           (103),
		.PKT_THREAD_ID_L           (103),
		.PKT_CACHE_H               (110),
		.PKT_CACHE_L               (107),
		.PKT_DATA_SIDEBAND_H       (92),
		.PKT_DATA_SIDEBAND_L       (92),
		.PKT_QOS_H                 (94),
		.PKT_QOS_L                 (94),
		.PKT_ADDR_SIDEBAND_H       (91),
		.PKT_ADDR_SIDEBAND_L       (91),
		.ST_DATA_W                 (113),
		.ST_CHANNEL_W              (12),
		.AV_BURSTCOUNT_W           (6),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (1),
		.BURSTWRAP_VALUE           (63),
		.CACHE_VALUE               (4'b0000)
	) com_nios_data_master_translator_avalon_universal_master_0_agent (
		.clk              (clk_clk),                                                                          //       clk.clk
		.reset            (rst_controller_reset_out_reset),                                                   // clk_reset.reset
		.av_address       (com_nios_data_master_translator_avalon_universal_master_0_address),                //        av.address
		.av_write         (com_nios_data_master_translator_avalon_universal_master_0_write),                  //          .write
		.av_read          (com_nios_data_master_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata     (com_nios_data_master_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata      (com_nios_data_master_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest   (com_nios_data_master_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid (com_nios_data_master_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable    (com_nios_data_master_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount    (com_nios_data_master_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess   (com_nios_data_master_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock          (com_nios_data_master_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid         (com_nios_data_master_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data          (com_nios_data_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket (com_nios_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket   (com_nios_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready         (com_nios_data_master_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid         (limiter_001_rsp_src_valid),                                                        //        rp.valid
		.rp_data          (limiter_001_rsp_src_data),                                                         //          .data
		.rp_channel       (limiter_001_rsp_src_channel),                                                      //          .channel
		.rp_startofpacket (limiter_001_rsp_src_startofpacket),                                                //          .startofpacket
		.rp_endofpacket   (limiter_001_rsp_src_endofpacket),                                                  //          .endofpacket
		.rp_ready         (limiter_001_rsp_src_ready)                                                         //          .ready
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (106),
		.PKT_PROTECTION_L          (104),
		.PKT_BEGIN_BURST           (93),
		.PKT_BURSTWRAP_H           (85),
		.PKT_BURSTWRAP_L           (80),
		.PKT_BURST_SIZE_H          (88),
		.PKT_BURST_SIZE_L          (86),
		.PKT_BURST_TYPE_H          (90),
		.PKT_BURST_TYPE_L          (89),
		.PKT_BYTE_CNT_H            (79),
		.PKT_BYTE_CNT_L            (74),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_TRANS_EXCLUSIVE       (73),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (98),
		.PKT_SRC_ID_L              (95),
		.PKT_DEST_ID_H             (102),
		.PKT_DEST_ID_L             (99),
		.PKT_THREAD_ID_H           (103),
		.PKT_THREAD_ID_L           (103),
		.PKT_CACHE_H               (110),
		.PKT_CACHE_L               (107),
		.PKT_DATA_SIDEBAND_H       (92),
		.PKT_DATA_SIDEBAND_L       (92),
		.PKT_QOS_H                 (94),
		.PKT_QOS_L                 (94),
		.PKT_ADDR_SIDEBAND_H       (91),
		.PKT_ADDR_SIDEBAND_L       (91),
		.ST_DATA_W                 (113),
		.ST_CHANNEL_W              (12),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (2),
		.BURSTWRAP_VALUE           (63),
		.CACHE_VALUE               (4'b0000)
	) carcontrol_nios_data_master_translator_avalon_universal_master_0_agent (
		.clk              (clk_clk),                                                                                 //       clk.clk
		.reset            (rst_controller_reset_out_reset),                                                          // clk_reset.reset
		.av_address       (carcontrol_nios_data_master_translator_avalon_universal_master_0_address),                //        av.address
		.av_write         (carcontrol_nios_data_master_translator_avalon_universal_master_0_write),                  //          .write
		.av_read          (carcontrol_nios_data_master_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata     (carcontrol_nios_data_master_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata      (carcontrol_nios_data_master_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest   (carcontrol_nios_data_master_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid (carcontrol_nios_data_master_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable    (carcontrol_nios_data_master_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount    (carcontrol_nios_data_master_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess   (carcontrol_nios_data_master_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock          (carcontrol_nios_data_master_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid         (carcontrol_nios_data_master_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data          (carcontrol_nios_data_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket (carcontrol_nios_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket   (carcontrol_nios_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready         (carcontrol_nios_data_master_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid         (rsp_xbar_mux_002_src_valid),                                                              //        rp.valid
		.rp_data          (rsp_xbar_mux_002_src_data),                                                               //          .data
		.rp_channel       (rsp_xbar_mux_002_src_channel),                                                            //          .channel
		.rp_startofpacket (rsp_xbar_mux_002_src_startofpacket),                                                      //          .startofpacket
		.rp_endofpacket   (rsp_xbar_mux_002_src_endofpacket),                                                        //          .endofpacket
		.rp_ready         (rsp_xbar_mux_002_src_ready)                                                               //          .ready
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (106),
		.PKT_PROTECTION_L          (104),
		.PKT_BEGIN_BURST           (93),
		.PKT_BURSTWRAP_H           (85),
		.PKT_BURSTWRAP_L           (80),
		.PKT_BURST_SIZE_H          (88),
		.PKT_BURST_SIZE_L          (86),
		.PKT_BURST_TYPE_H          (90),
		.PKT_BURST_TYPE_L          (89),
		.PKT_BYTE_CNT_H            (79),
		.PKT_BYTE_CNT_L            (74),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_TRANS_EXCLUSIVE       (73),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (98),
		.PKT_SRC_ID_L              (95),
		.PKT_DEST_ID_H             (102),
		.PKT_DEST_ID_L             (99),
		.PKT_THREAD_ID_H           (103),
		.PKT_THREAD_ID_L           (103),
		.PKT_CACHE_H               (110),
		.PKT_CACHE_L               (107),
		.PKT_DATA_SIDEBAND_H       (92),
		.PKT_DATA_SIDEBAND_L       (92),
		.PKT_QOS_H                 (94),
		.PKT_QOS_L                 (94),
		.PKT_ADDR_SIDEBAND_H       (91),
		.PKT_ADDR_SIDEBAND_L       (91),
		.ST_DATA_W                 (113),
		.ST_CHANNEL_W              (12),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (3),
		.BURSTWRAP_VALUE           (3),
		.CACHE_VALUE               (4'b0000)
	) carcontrol_nios_instruction_master_translator_avalon_universal_master_0_agent (
		.clk              (clk_clk),                                                                                        //       clk.clk
		.reset            (rst_controller_reset_out_reset),                                                                 // clk_reset.reset
		.av_address       (carcontrol_nios_instruction_master_translator_avalon_universal_master_0_address),                //        av.address
		.av_write         (carcontrol_nios_instruction_master_translator_avalon_universal_master_0_write),                  //          .write
		.av_read          (carcontrol_nios_instruction_master_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata     (carcontrol_nios_instruction_master_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata      (carcontrol_nios_instruction_master_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest   (carcontrol_nios_instruction_master_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid (carcontrol_nios_instruction_master_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable    (carcontrol_nios_instruction_master_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount    (carcontrol_nios_instruction_master_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess   (carcontrol_nios_instruction_master_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock          (carcontrol_nios_instruction_master_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid         (carcontrol_nios_instruction_master_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data          (carcontrol_nios_instruction_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket (carcontrol_nios_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket   (carcontrol_nios_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready         (carcontrol_nios_instruction_master_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid         (limiter_002_rsp_src_valid),                                                                      //        rp.valid
		.rp_data          (limiter_002_rsp_src_data),                                                                       //          .data
		.rp_channel       (limiter_002_rsp_src_channel),                                                                    //          .channel
		.rp_startofpacket (limiter_002_rsp_src_startofpacket),                                                              //          .startofpacket
		.rp_endofpacket   (limiter_002_rsp_src_endofpacket),                                                                //          .endofpacket
		.rp_ready         (limiter_002_rsp_src_ready)                                                                       //          .ready
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (106),
		.PKT_PROTECTION_L          (104),
		.PKT_BEGIN_BURST           (93),
		.PKT_BURSTWRAP_H           (85),
		.PKT_BURSTWRAP_L           (80),
		.PKT_BURST_SIZE_H          (88),
		.PKT_BURST_SIZE_L          (86),
		.PKT_BURST_TYPE_H          (90),
		.PKT_BURST_TYPE_L          (89),
		.PKT_BYTE_CNT_H            (79),
		.PKT_BYTE_CNT_L            (74),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_TRANS_EXCLUSIVE       (73),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (98),
		.PKT_SRC_ID_L              (95),
		.PKT_DEST_ID_H             (102),
		.PKT_DEST_ID_L             (99),
		.PKT_THREAD_ID_H           (103),
		.PKT_THREAD_ID_L           (103),
		.PKT_CACHE_H               (110),
		.PKT_CACHE_L               (107),
		.PKT_DATA_SIDEBAND_H       (92),
		.PKT_DATA_SIDEBAND_L       (92),
		.PKT_QOS_H                 (94),
		.PKT_QOS_L                 (94),
		.PKT_ADDR_SIDEBAND_H       (91),
		.PKT_ADDR_SIDEBAND_L       (91),
		.ST_DATA_W                 (113),
		.ST_CHANNEL_W              (12),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (4),
		.BURSTWRAP_VALUE           (63),
		.CACHE_VALUE               (4'b0000)
	) ethernet_subsystem_sgdma_rx_m_write_translator_avalon_universal_master_0_agent (
		.clk              (clk_clk),                                                                                         //       clk.clk
		.reset            (rst_controller_002_reset_out_reset),                                                              // clk_reset.reset
		.av_address       (ethernet_subsystem_sgdma_rx_m_write_translator_avalon_universal_master_0_address),                //        av.address
		.av_write         (ethernet_subsystem_sgdma_rx_m_write_translator_avalon_universal_master_0_write),                  //          .write
		.av_read          (ethernet_subsystem_sgdma_rx_m_write_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata     (ethernet_subsystem_sgdma_rx_m_write_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata      (ethernet_subsystem_sgdma_rx_m_write_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest   (ethernet_subsystem_sgdma_rx_m_write_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid (ethernet_subsystem_sgdma_rx_m_write_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable    (ethernet_subsystem_sgdma_rx_m_write_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount    (ethernet_subsystem_sgdma_rx_m_write_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess   (ethernet_subsystem_sgdma_rx_m_write_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock          (ethernet_subsystem_sgdma_rx_m_write_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid         (ethernet_subsystem_sgdma_rx_m_write_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data          (ethernet_subsystem_sgdma_rx_m_write_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket (ethernet_subsystem_sgdma_rx_m_write_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket   (ethernet_subsystem_sgdma_rx_m_write_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready         (ethernet_subsystem_sgdma_rx_m_write_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid         (rsp_xbar_demux_001_src2_valid),                                                                   //        rp.valid
		.rp_data          (rsp_xbar_demux_001_src2_data),                                                                    //          .data
		.rp_channel       (rsp_xbar_demux_001_src2_channel),                                                                 //          .channel
		.rp_startofpacket (rsp_xbar_demux_001_src2_startofpacket),                                                           //          .startofpacket
		.rp_endofpacket   (rsp_xbar_demux_001_src2_endofpacket),                                                             //          .endofpacket
		.rp_ready         (rsp_xbar_demux_001_src2_ready)                                                                    //          .ready
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (106),
		.PKT_PROTECTION_L          (104),
		.PKT_BEGIN_BURST           (93),
		.PKT_BURSTWRAP_H           (85),
		.PKT_BURSTWRAP_L           (80),
		.PKT_BURST_SIZE_H          (88),
		.PKT_BURST_SIZE_L          (86),
		.PKT_BURST_TYPE_H          (90),
		.PKT_BURST_TYPE_L          (89),
		.PKT_BYTE_CNT_H            (79),
		.PKT_BYTE_CNT_L            (74),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_TRANS_EXCLUSIVE       (73),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (98),
		.PKT_SRC_ID_L              (95),
		.PKT_DEST_ID_H             (102),
		.PKT_DEST_ID_L             (99),
		.PKT_THREAD_ID_H           (103),
		.PKT_THREAD_ID_L           (103),
		.PKT_CACHE_H               (110),
		.PKT_CACHE_L               (107),
		.PKT_DATA_SIDEBAND_H       (92),
		.PKT_DATA_SIDEBAND_L       (92),
		.PKT_QOS_H                 (94),
		.PKT_QOS_L                 (94),
		.PKT_ADDR_SIDEBAND_H       (91),
		.PKT_ADDR_SIDEBAND_L       (91),
		.ST_DATA_W                 (113),
		.ST_CHANNEL_W              (12),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (5),
		.BURSTWRAP_VALUE           (63),
		.CACHE_VALUE               (4'b0000)
	) ethernet_subsystem_sgdma_tx_m_read_translator_avalon_universal_master_0_agent (
		.clk              (clk_clk),                                                                                        //       clk.clk
		.reset            (rst_controller_002_reset_out_reset),                                                             // clk_reset.reset
		.av_address       (ethernet_subsystem_sgdma_tx_m_read_translator_avalon_universal_master_0_address),                //        av.address
		.av_write         (ethernet_subsystem_sgdma_tx_m_read_translator_avalon_universal_master_0_write),                  //          .write
		.av_read          (ethernet_subsystem_sgdma_tx_m_read_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata     (ethernet_subsystem_sgdma_tx_m_read_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata      (ethernet_subsystem_sgdma_tx_m_read_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest   (ethernet_subsystem_sgdma_tx_m_read_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid (ethernet_subsystem_sgdma_tx_m_read_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable    (ethernet_subsystem_sgdma_tx_m_read_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount    (ethernet_subsystem_sgdma_tx_m_read_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess   (ethernet_subsystem_sgdma_tx_m_read_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock          (ethernet_subsystem_sgdma_tx_m_read_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid         (ethernet_subsystem_sgdma_tx_m_read_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data          (ethernet_subsystem_sgdma_tx_m_read_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket (ethernet_subsystem_sgdma_tx_m_read_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket   (ethernet_subsystem_sgdma_tx_m_read_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready         (ethernet_subsystem_sgdma_tx_m_read_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid         (rsp_xbar_demux_001_src3_valid),                                                                  //        rp.valid
		.rp_data          (rsp_xbar_demux_001_src3_data),                                                                   //          .data
		.rp_channel       (rsp_xbar_demux_001_src3_channel),                                                                //          .channel
		.rp_startofpacket (rsp_xbar_demux_001_src3_startofpacket),                                                          //          .startofpacket
		.rp_endofpacket   (rsp_xbar_demux_001_src3_endofpacket),                                                            //          .endofpacket
		.rp_ready         (rsp_xbar_demux_001_src3_ready)                                                                   //          .ready
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (93),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (98),
		.PKT_SRC_ID_L              (95),
		.PKT_DEST_ID_H             (102),
		.PKT_DEST_ID_L             (99),
		.PKT_BURSTWRAP_H           (85),
		.PKT_BURSTWRAP_L           (80),
		.PKT_BYTE_CNT_H            (79),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (106),
		.PKT_PROTECTION_L          (104),
		.PKT_RESPONSE_STATUS_H     (112),
		.PKT_RESPONSE_STATUS_L     (111),
		.PKT_BURST_SIZE_H          (88),
		.PKT_BURST_SIZE_L          (86),
		.ST_CHANNEL_W              (12),
		.ST_DATA_W                 (113),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) com_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                         //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                                  //       clk_reset.reset
		.m0_address              (com_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (com_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (com_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (com_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (com_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (com_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (com_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (com_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (com_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (com_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (com_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (com_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (com_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (com_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (com_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (com_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (burst_adapter_source0_ready),                                                                     //              cp.ready
		.cp_valid                (burst_adapter_source0_valid),                                                                     //                .valid
		.cp_data                 (burst_adapter_source0_data),                                                                      //                .data
		.cp_startofpacket        (burst_adapter_source0_startofpacket),                                                             //                .startofpacket
		.cp_endofpacket          (burst_adapter_source0_endofpacket),                                                               //                .endofpacket
		.cp_channel              (burst_adapter_source0_channel),                                                                   //                .channel
		.rf_sink_ready           (com_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (com_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (com_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (com_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (com_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (com_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (com_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (com_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (com_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (com_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (com_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (com_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (com_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (com_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (com_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (com_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (114),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) com_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                         //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                                  // clk_reset.reset
		.in_data           (com_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (com_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (com_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (com_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (com_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (com_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (com_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (com_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (com_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (com_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                           // (terminated)
		.csr_read          (1'b0),                                                                                            // (terminated)
		.csr_write         (1'b0),                                                                                            // (terminated)
		.csr_readdata      (),                                                                                                // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                            // (terminated)
		.almost_full_data  (),                                                                                                // (terminated)
		.almost_empty_data (),                                                                                                // (terminated)
		.in_empty          (1'b0),                                                                                            // (terminated)
		.out_empty         (),                                                                                                // (terminated)
		.in_error          (1'b0),                                                                                            // (terminated)
		.out_error         (),                                                                                                // (terminated)
		.in_channel        (1'b0),                                                                                            // (terminated)
		.out_channel       ()                                                                                                 // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (93),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (98),
		.PKT_SRC_ID_L              (95),
		.PKT_DEST_ID_H             (102),
		.PKT_DEST_ID_L             (99),
		.PKT_BURSTWRAP_H           (85),
		.PKT_BURSTWRAP_L           (80),
		.PKT_BYTE_CNT_H            (79),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (106),
		.PKT_PROTECTION_L          (104),
		.PKT_RESPONSE_STATUS_H     (112),
		.PKT_RESPONSE_STATUS_L     (111),
		.PKT_BURST_SIZE_H          (88),
		.PKT_BURST_SIZE_L          (86),
		.ST_CHANNEL_W              (12),
		.ST_DATA_W                 (113),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) com_memory_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                            //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                     //       clk_reset.reset
		.m0_address              (com_memory_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (com_memory_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (com_memory_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (com_memory_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (com_memory_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (com_memory_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (com_memory_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (com_memory_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (com_memory_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (com_memory_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (com_memory_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (com_memory_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (com_memory_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (com_memory_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (com_memory_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (com_memory_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (burst_adapter_001_source0_ready),                                                    //              cp.ready
		.cp_valid                (burst_adapter_001_source0_valid),                                                    //                .valid
		.cp_data                 (burst_adapter_001_source0_data),                                                     //                .data
		.cp_startofpacket        (burst_adapter_001_source0_startofpacket),                                            //                .startofpacket
		.cp_endofpacket          (burst_adapter_001_source0_endofpacket),                                              //                .endofpacket
		.cp_channel              (burst_adapter_001_source0_channel),                                                  //                .channel
		.rf_sink_ready           (com_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (com_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (com_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (com_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (com_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (com_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (com_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (com_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (com_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (com_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (com_memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (com_memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (com_memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (com_memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (com_memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (com_memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (114),
		.FIFO_DEPTH          (8),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) com_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                            //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                     // clk_reset.reset
		.in_data           (com_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (com_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (com_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (com_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (com_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (com_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (com_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (com_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (com_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (com_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                              // (terminated)
		.csr_read          (1'b0),                                                                               // (terminated)
		.csr_write         (1'b0),                                                                               // (terminated)
		.csr_readdata      (),                                                                                   // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                               // (terminated)
		.almost_full_data  (),                                                                                   // (terminated)
		.almost_empty_data (),                                                                                   // (terminated)
		.in_empty          (1'b0),                                                                               // (terminated)
		.out_empty         (),                                                                                   // (terminated)
		.in_error          (1'b0),                                                                               // (terminated)
		.out_error         (),                                                                                   // (terminated)
		.in_channel        (1'b0),                                                                               // (terminated)
		.out_channel       ()                                                                                    // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (93),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (98),
		.PKT_SRC_ID_L              (95),
		.PKT_DEST_ID_H             (102),
		.PKT_DEST_ID_L             (99),
		.PKT_BURSTWRAP_H           (85),
		.PKT_BURSTWRAP_L           (80),
		.PKT_BYTE_CNT_H            (79),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (106),
		.PKT_PROTECTION_L          (104),
		.PKT_RESPONSE_STATUS_H     (112),
		.PKT_RESPONSE_STATUS_L     (111),
		.PKT_BURST_SIZE_H          (88),
		.PKT_BURST_SIZE_L          (86),
		.ST_CHANNEL_W              (12),
		.ST_DATA_W                 (113),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) jtaguart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                           //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                                //       clk_reset.reset
		.m0_address              (jtaguart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (jtaguart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (jtaguart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (jtaguart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (jtaguart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (jtaguart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (jtaguart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (jtaguart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (jtaguart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (jtaguart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (jtaguart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (jtaguart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (jtaguart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (jtaguart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (jtaguart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (jtaguart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (burst_adapter_002_source0_ready),                                                                   //              cp.ready
		.cp_valid                (burst_adapter_002_source0_valid),                                                                   //                .valid
		.cp_data                 (burst_adapter_002_source0_data),                                                                    //                .data
		.cp_startofpacket        (burst_adapter_002_source0_startofpacket),                                                           //                .startofpacket
		.cp_endofpacket          (burst_adapter_002_source0_endofpacket),                                                             //                .endofpacket
		.cp_channel              (burst_adapter_002_source0_channel),                                                                 //                .channel
		.rf_sink_ready           (jtaguart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (jtaguart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (jtaguart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (jtaguart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (jtaguart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (jtaguart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (jtaguart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (jtaguart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (jtaguart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (jtaguart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (jtaguart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (jtaguart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (jtaguart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (jtaguart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (jtaguart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (jtaguart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (114),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) jtaguart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                           //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                                // clk_reset.reset
		.in_data           (jtaguart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (jtaguart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (jtaguart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (jtaguart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (jtaguart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (jtaguart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (jtaguart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (jtaguart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (jtaguart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (jtaguart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                             // (terminated)
		.csr_read          (1'b0),                                                                                              // (terminated)
		.csr_write         (1'b0),                                                                                              // (terminated)
		.csr_readdata      (),                                                                                                  // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                              // (terminated)
		.almost_full_data  (),                                                                                                  // (terminated)
		.almost_empty_data (),                                                                                                  // (terminated)
		.in_empty          (1'b0),                                                                                              // (terminated)
		.out_empty         (),                                                                                                  // (terminated)
		.in_error          (1'b0),                                                                                              // (terminated)
		.out_error         (),                                                                                                  // (terminated)
		.in_channel        (1'b0),                                                                                              // (terminated)
		.out_channel       ()                                                                                                   // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (93),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (98),
		.PKT_SRC_ID_L              (95),
		.PKT_DEST_ID_H             (102),
		.PKT_DEST_ID_L             (99),
		.PKT_BURSTWRAP_H           (85),
		.PKT_BURSTWRAP_L           (80),
		.PKT_BYTE_CNT_H            (79),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (106),
		.PKT_PROTECTION_L          (104),
		.PKT_RESPONSE_STATUS_H     (112),
		.PKT_RESPONSE_STATUS_L     (111),
		.PKT_BURST_SIZE_H          (88),
		.PKT_BURST_SIZE_L          (86),
		.ST_CHANNEL_W              (12),
		.ST_DATA_W                 (113),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) shared_memory_mutex_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                     //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                              //       clk_reset.reset
		.m0_address              (shared_memory_mutex_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (shared_memory_mutex_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (shared_memory_mutex_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (shared_memory_mutex_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (shared_memory_mutex_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (shared_memory_mutex_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (shared_memory_mutex_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (shared_memory_mutex_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (shared_memory_mutex_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (shared_memory_mutex_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (shared_memory_mutex_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (shared_memory_mutex_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (shared_memory_mutex_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (shared_memory_mutex_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (shared_memory_mutex_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (shared_memory_mutex_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (burst_adapter_003_source0_ready),                                                             //              cp.ready
		.cp_valid                (burst_adapter_003_source0_valid),                                                             //                .valid
		.cp_data                 (burst_adapter_003_source0_data),                                                              //                .data
		.cp_startofpacket        (burst_adapter_003_source0_startofpacket),                                                     //                .startofpacket
		.cp_endofpacket          (burst_adapter_003_source0_endofpacket),                                                       //                .endofpacket
		.cp_channel              (burst_adapter_003_source0_channel),                                                           //                .channel
		.rf_sink_ready           (shared_memory_mutex_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (shared_memory_mutex_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (shared_memory_mutex_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (shared_memory_mutex_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (shared_memory_mutex_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (shared_memory_mutex_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (shared_memory_mutex_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (shared_memory_mutex_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (shared_memory_mutex_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (shared_memory_mutex_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (shared_memory_mutex_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (shared_memory_mutex_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (shared_memory_mutex_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (shared_memory_mutex_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (shared_memory_mutex_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (shared_memory_mutex_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (114),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) shared_memory_mutex_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                     //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                              // clk_reset.reset
		.in_data           (shared_memory_mutex_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (shared_memory_mutex_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (shared_memory_mutex_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (shared_memory_mutex_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (shared_memory_mutex_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (shared_memory_mutex_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (shared_memory_mutex_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (shared_memory_mutex_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (shared_memory_mutex_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (shared_memory_mutex_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                       // (terminated)
		.csr_read          (1'b0),                                                                                        // (terminated)
		.csr_write         (1'b0),                                                                                        // (terminated)
		.csr_readdata      (),                                                                                            // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                        // (terminated)
		.almost_full_data  (),                                                                                            // (terminated)
		.almost_empty_data (),                                                                                            // (terminated)
		.in_empty          (1'b0),                                                                                        // (terminated)
		.out_empty         (),                                                                                            // (terminated)
		.in_error          (1'b0),                                                                                        // (terminated)
		.out_error         (),                                                                                            // (terminated)
		.in_channel        (1'b0),                                                                                        // (terminated)
		.out_channel       ()                                                                                             // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (93),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (98),
		.PKT_SRC_ID_L              (95),
		.PKT_DEST_ID_H             (102),
		.PKT_DEST_ID_L             (99),
		.PKT_BURSTWRAP_H           (85),
		.PKT_BURSTWRAP_L           (80),
		.PKT_BYTE_CNT_H            (79),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (106),
		.PKT_PROTECTION_L          (104),
		.PKT_RESPONSE_STATUS_H     (112),
		.PKT_RESPONSE_STATUS_L     (111),
		.PKT_BURST_SIZE_H          (88),
		.PKT_BURST_SIZE_L          (86),
		.ST_CHANNEL_W              (12),
		.ST_DATA_W                 (113),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) com_timer_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                           //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                    //       clk_reset.reset
		.m0_address              (com_timer_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (com_timer_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (com_timer_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (com_timer_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (com_timer_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (com_timer_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (com_timer_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (com_timer_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (com_timer_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (com_timer_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (com_timer_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (com_timer_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (com_timer_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (com_timer_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (com_timer_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (com_timer_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (burst_adapter_004_source0_ready),                                                   //              cp.ready
		.cp_valid                (burst_adapter_004_source0_valid),                                                   //                .valid
		.cp_data                 (burst_adapter_004_source0_data),                                                    //                .data
		.cp_startofpacket        (burst_adapter_004_source0_startofpacket),                                           //                .startofpacket
		.cp_endofpacket          (burst_adapter_004_source0_endofpacket),                                             //                .endofpacket
		.cp_channel              (burst_adapter_004_source0_channel),                                                 //                .channel
		.rf_sink_ready           (com_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (com_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (com_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (com_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (com_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (com_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (com_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (com_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (com_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (com_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (com_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (com_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (com_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (com_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (com_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (com_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (114),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) com_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                           //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                    // clk_reset.reset
		.in_data           (com_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (com_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (com_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (com_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (com_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (com_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (com_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (com_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (com_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (com_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                             // (terminated)
		.csr_read          (1'b0),                                                                              // (terminated)
		.csr_write         (1'b0),                                                                              // (terminated)
		.csr_readdata      (),                                                                                  // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                              // (terminated)
		.almost_full_data  (),                                                                                  // (terminated)
		.almost_empty_data (),                                                                                  // (terminated)
		.in_empty          (1'b0),                                                                              // (terminated)
		.out_empty         (),                                                                                  // (terminated)
		.in_error          (1'b0),                                                                              // (terminated)
		.out_error         (),                                                                                  // (terminated)
		.in_channel        (1'b0),                                                                              // (terminated)
		.out_channel       ()                                                                                   // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (93),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (98),
		.PKT_SRC_ID_L              (95),
		.PKT_DEST_ID_H             (102),
		.PKT_DEST_ID_L             (99),
		.PKT_BURSTWRAP_H           (85),
		.PKT_BURSTWRAP_L           (80),
		.PKT_BYTE_CNT_H            (79),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (106),
		.PKT_PROTECTION_L          (104),
		.PKT_RESPONSE_STATUS_H     (112),
		.PKT_RESPONSE_STATUS_L     (111),
		.PKT_BURST_SIZE_H          (88),
		.PKT_BURST_SIZE_L          (86),
		.ST_CHANNEL_W              (12),
		.ST_DATA_W                 (113),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) ethernet_subsystem_ethernet_bridge_s0_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                                    //             clk.clk
		.reset                   (rst_controller_002_reset_out_reset),                                                                         //       clk_reset.reset
		.m0_address              (ethernet_subsystem_ethernet_bridge_s0_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (ethernet_subsystem_ethernet_bridge_s0_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (ethernet_subsystem_ethernet_bridge_s0_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (ethernet_subsystem_ethernet_bridge_s0_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (ethernet_subsystem_ethernet_bridge_s0_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (ethernet_subsystem_ethernet_bridge_s0_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (ethernet_subsystem_ethernet_bridge_s0_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (ethernet_subsystem_ethernet_bridge_s0_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (ethernet_subsystem_ethernet_bridge_s0_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (ethernet_subsystem_ethernet_bridge_s0_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (ethernet_subsystem_ethernet_bridge_s0_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (ethernet_subsystem_ethernet_bridge_s0_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (ethernet_subsystem_ethernet_bridge_s0_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (ethernet_subsystem_ethernet_bridge_s0_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (ethernet_subsystem_ethernet_bridge_s0_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (ethernet_subsystem_ethernet_bridge_s0_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (burst_adapter_005_source0_ready),                                                                            //              cp.ready
		.cp_valid                (burst_adapter_005_source0_valid),                                                                            //                .valid
		.cp_data                 (burst_adapter_005_source0_data),                                                                             //                .data
		.cp_startofpacket        (burst_adapter_005_source0_startofpacket),                                                                    //                .startofpacket
		.cp_endofpacket          (burst_adapter_005_source0_endofpacket),                                                                      //                .endofpacket
		.cp_channel              (burst_adapter_005_source0_channel),                                                                          //                .channel
		.rf_sink_ready           (ethernet_subsystem_ethernet_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (ethernet_subsystem_ethernet_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (ethernet_subsystem_ethernet_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (ethernet_subsystem_ethernet_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (ethernet_subsystem_ethernet_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (ethernet_subsystem_ethernet_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (ethernet_subsystem_ethernet_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (ethernet_subsystem_ethernet_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (ethernet_subsystem_ethernet_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (ethernet_subsystem_ethernet_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (ethernet_subsystem_ethernet_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (ethernet_subsystem_ethernet_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (ethernet_subsystem_ethernet_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (ethernet_subsystem_ethernet_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (ethernet_subsystem_ethernet_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (ethernet_subsystem_ethernet_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (114),
		.FIFO_DEPTH          (5),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) ethernet_subsystem_ethernet_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                                    //       clk.clk
		.reset             (rst_controller_002_reset_out_reset),                                                                         // clk_reset.reset
		.in_data           (ethernet_subsystem_ethernet_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (ethernet_subsystem_ethernet_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (ethernet_subsystem_ethernet_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (ethernet_subsystem_ethernet_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (ethernet_subsystem_ethernet_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (ethernet_subsystem_ethernet_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (ethernet_subsystem_ethernet_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (ethernet_subsystem_ethernet_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (ethernet_subsystem_ethernet_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (ethernet_subsystem_ethernet_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                                      // (terminated)
		.csr_read          (1'b0),                                                                                                       // (terminated)
		.csr_write         (1'b0),                                                                                                       // (terminated)
		.csr_readdata      (),                                                                                                           // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                                       // (terminated)
		.almost_full_data  (),                                                                                                           // (terminated)
		.almost_empty_data (),                                                                                                           // (terminated)
		.in_empty          (1'b0),                                                                                                       // (terminated)
		.out_empty         (),                                                                                                           // (terminated)
		.in_error          (1'b0),                                                                                                       // (terminated)
		.out_error         (),                                                                                                           // (terminated)
		.in_channel        (1'b0),                                                                                                       // (terminated)
		.out_channel       ()                                                                                                            // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (93),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (98),
		.PKT_SRC_ID_L              (95),
		.PKT_DEST_ID_H             (102),
		.PKT_DEST_ID_L             (99),
		.PKT_BURSTWRAP_H           (85),
		.PKT_BURSTWRAP_L           (80),
		.PKT_BYTE_CNT_H            (79),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (106),
		.PKT_PROTECTION_L          (104),
		.PKT_RESPONSE_STATUS_H     (112),
		.PKT_RESPONSE_STATUS_L     (111),
		.PKT_BURST_SIZE_H          (88),
		.PKT_BURST_SIZE_L          (86),
		.ST_CHANNEL_W              (12),
		.ST_DATA_W                 (113),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) ethernet_subsystem_descriptor_memory_s2_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                                      //             clk.clk
		.reset                   (rst_controller_002_reset_out_reset),                                                                           //       clk_reset.reset
		.m0_address              (ethernet_subsystem_descriptor_memory_s2_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (ethernet_subsystem_descriptor_memory_s2_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (ethernet_subsystem_descriptor_memory_s2_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (ethernet_subsystem_descriptor_memory_s2_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (ethernet_subsystem_descriptor_memory_s2_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (ethernet_subsystem_descriptor_memory_s2_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (ethernet_subsystem_descriptor_memory_s2_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (ethernet_subsystem_descriptor_memory_s2_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (ethernet_subsystem_descriptor_memory_s2_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (ethernet_subsystem_descriptor_memory_s2_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (ethernet_subsystem_descriptor_memory_s2_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (ethernet_subsystem_descriptor_memory_s2_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (ethernet_subsystem_descriptor_memory_s2_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (ethernet_subsystem_descriptor_memory_s2_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (ethernet_subsystem_descriptor_memory_s2_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (ethernet_subsystem_descriptor_memory_s2_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (burst_adapter_006_source0_ready),                                                                              //              cp.ready
		.cp_valid                (burst_adapter_006_source0_valid),                                                                              //                .valid
		.cp_data                 (burst_adapter_006_source0_data),                                                                               //                .data
		.cp_startofpacket        (burst_adapter_006_source0_startofpacket),                                                                      //                .startofpacket
		.cp_endofpacket          (burst_adapter_006_source0_endofpacket),                                                                        //                .endofpacket
		.cp_channel              (burst_adapter_006_source0_channel),                                                                            //                .channel
		.rf_sink_ready           (ethernet_subsystem_descriptor_memory_s2_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (ethernet_subsystem_descriptor_memory_s2_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (ethernet_subsystem_descriptor_memory_s2_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (ethernet_subsystem_descriptor_memory_s2_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (ethernet_subsystem_descriptor_memory_s2_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (ethernet_subsystem_descriptor_memory_s2_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (ethernet_subsystem_descriptor_memory_s2_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (ethernet_subsystem_descriptor_memory_s2_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (ethernet_subsystem_descriptor_memory_s2_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (ethernet_subsystem_descriptor_memory_s2_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (ethernet_subsystem_descriptor_memory_s2_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (ethernet_subsystem_descriptor_memory_s2_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (ethernet_subsystem_descriptor_memory_s2_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (ethernet_subsystem_descriptor_memory_s2_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (ethernet_subsystem_descriptor_memory_s2_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (ethernet_subsystem_descriptor_memory_s2_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (114),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) ethernet_subsystem_descriptor_memory_s2_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                                      //       clk.clk
		.reset             (rst_controller_002_reset_out_reset),                                                                           // clk_reset.reset
		.in_data           (ethernet_subsystem_descriptor_memory_s2_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (ethernet_subsystem_descriptor_memory_s2_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (ethernet_subsystem_descriptor_memory_s2_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (ethernet_subsystem_descriptor_memory_s2_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (ethernet_subsystem_descriptor_memory_s2_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (ethernet_subsystem_descriptor_memory_s2_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (ethernet_subsystem_descriptor_memory_s2_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (ethernet_subsystem_descriptor_memory_s2_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (ethernet_subsystem_descriptor_memory_s2_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (ethernet_subsystem_descriptor_memory_s2_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                                        // (terminated)
		.csr_read          (1'b0),                                                                                                         // (terminated)
		.csr_write         (1'b0),                                                                                                         // (terminated)
		.csr_readdata      (),                                                                                                             // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                                         // (terminated)
		.almost_full_data  (),                                                                                                             // (terminated)
		.almost_empty_data (),                                                                                                             // (terminated)
		.in_empty          (1'b0),                                                                                                         // (terminated)
		.out_empty         (),                                                                                                             // (terminated)
		.in_error          (1'b0),                                                                                                         // (terminated)
		.out_error         (),                                                                                                             // (terminated)
		.in_channel        (1'b0),                                                                                                         // (terminated)
		.out_channel       ()                                                                                                              // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (93),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (98),
		.PKT_SRC_ID_L              (95),
		.PKT_DEST_ID_H             (102),
		.PKT_DEST_ID_L             (99),
		.PKT_BURSTWRAP_H           (85),
		.PKT_BURSTWRAP_L           (80),
		.PKT_BYTE_CNT_H            (79),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (106),
		.PKT_PROTECTION_L          (104),
		.PKT_RESPONSE_STATUS_H     (112),
		.PKT_RESPONSE_STATUS_L     (111),
		.PKT_BURST_SIZE_H          (88),
		.PKT_BURST_SIZE_L          (86),
		.ST_CHANNEL_W              (12),
		.ST_DATA_W                 (113),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) prio_arbiter_0_s0_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                         //       clk_reset.reset
		.m0_address              (prio_arbiter_0_s0_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (prio_arbiter_0_s0_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (prio_arbiter_0_s0_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (prio_arbiter_0_s0_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (prio_arbiter_0_s0_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (prio_arbiter_0_s0_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (prio_arbiter_0_s0_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (prio_arbiter_0_s0_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (prio_arbiter_0_s0_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (prio_arbiter_0_s0_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (prio_arbiter_0_s0_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (prio_arbiter_0_s0_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (prio_arbiter_0_s0_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (prio_arbiter_0_s0_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (prio_arbiter_0_s0_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (prio_arbiter_0_s0_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (burst_adapter_007_source0_ready),                                                        //              cp.ready
		.cp_valid                (burst_adapter_007_source0_valid),                                                        //                .valid
		.cp_data                 (burst_adapter_007_source0_data),                                                         //                .data
		.cp_startofpacket        (burst_adapter_007_source0_startofpacket),                                                //                .startofpacket
		.cp_endofpacket          (burst_adapter_007_source0_endofpacket),                                                  //                .endofpacket
		.cp_channel              (burst_adapter_007_source0_channel),                                                      //                .channel
		.rf_sink_ready           (prio_arbiter_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (prio_arbiter_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (prio_arbiter_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (prio_arbiter_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (prio_arbiter_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (prio_arbiter_0_s0_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (prio_arbiter_0_s0_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (prio_arbiter_0_s0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (prio_arbiter_0_s0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (prio_arbiter_0_s0_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (prio_arbiter_0_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (prio_arbiter_0_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (prio_arbiter_0_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (prio_arbiter_0_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (prio_arbiter_0_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (prio_arbiter_0_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (114),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) prio_arbiter_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                         // clk_reset.reset
		.in_data           (prio_arbiter_0_s0_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (prio_arbiter_0_s0_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (prio_arbiter_0_s0_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (prio_arbiter_0_s0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (prio_arbiter_0_s0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (prio_arbiter_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (prio_arbiter_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (prio_arbiter_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (prio_arbiter_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (prio_arbiter_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                  // (terminated)
		.csr_read          (1'b0),                                                                                   // (terminated)
		.csr_write         (1'b0),                                                                                   // (terminated)
		.csr_readdata      (),                                                                                       // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                   // (terminated)
		.almost_full_data  (),                                                                                       // (terminated)
		.almost_empty_data (),                                                                                       // (terminated)
		.in_empty          (1'b0),                                                                                   // (terminated)
		.out_empty         (),                                                                                       // (terminated)
		.in_error          (1'b0),                                                                                   // (terminated)
		.out_error         (),                                                                                       // (terminated)
		.in_channel        (1'b0),                                                                                   // (terminated)
		.out_channel       ()                                                                                        // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (93),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (98),
		.PKT_SRC_ID_L              (95),
		.PKT_DEST_ID_H             (102),
		.PKT_DEST_ID_L             (99),
		.PKT_BURSTWRAP_H           (85),
		.PKT_BURSTWRAP_L           (80),
		.PKT_BYTE_CNT_H            (79),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (106),
		.PKT_PROTECTION_L          (104),
		.PKT_RESPONSE_STATUS_H     (112),
		.PKT_RESPONSE_STATUS_L     (111),
		.PKT_BURST_SIZE_H          (88),
		.PKT_BURST_SIZE_L          (86),
		.ST_CHANNEL_W              (12),
		.ST_DATA_W                 (113),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) carcontrol_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                                //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                                         //       clk_reset.reset
		.m0_address              (carcontrol_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (carcontrol_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (carcontrol_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (carcontrol_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (carcontrol_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (carcontrol_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (carcontrol_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (carcontrol_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (carcontrol_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (carcontrol_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (carcontrol_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (carcontrol_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (carcontrol_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (carcontrol_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (carcontrol_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (carcontrol_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_008_src_ready),                                                                             //              cp.ready
		.cp_valid                (cmd_xbar_mux_008_src_valid),                                                                             //                .valid
		.cp_data                 (cmd_xbar_mux_008_src_data),                                                                              //                .data
		.cp_startofpacket        (cmd_xbar_mux_008_src_startofpacket),                                                                     //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_008_src_endofpacket),                                                                       //                .endofpacket
		.cp_channel              (cmd_xbar_mux_008_src_channel),                                                                           //                .channel
		.rf_sink_ready           (carcontrol_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (carcontrol_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (carcontrol_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (carcontrol_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (carcontrol_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (carcontrol_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (carcontrol_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (carcontrol_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (carcontrol_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (carcontrol_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (carcontrol_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (carcontrol_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (carcontrol_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (carcontrol_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (carcontrol_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (carcontrol_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (114),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) carcontrol_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                                //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                                         // clk_reset.reset
		.in_data           (carcontrol_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (carcontrol_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (carcontrol_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (carcontrol_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (carcontrol_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (carcontrol_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (carcontrol_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (carcontrol_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (carcontrol_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (carcontrol_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                                  // (terminated)
		.csr_read          (1'b0),                                                                                                   // (terminated)
		.csr_write         (1'b0),                                                                                                   // (terminated)
		.csr_readdata      (),                                                                                                       // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                                   // (terminated)
		.almost_full_data  (),                                                                                                       // (terminated)
		.almost_empty_data (),                                                                                                       // (terminated)
		.in_empty          (1'b0),                                                                                                   // (terminated)
		.out_empty         (),                                                                                                       // (terminated)
		.in_error          (1'b0),                                                                                                   // (terminated)
		.out_error         (),                                                                                                       // (terminated)
		.in_channel        (1'b0),                                                                                                   // (terminated)
		.out_channel       ()                                                                                                        // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (93),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (98),
		.PKT_SRC_ID_L              (95),
		.PKT_DEST_ID_H             (102),
		.PKT_DEST_ID_L             (99),
		.PKT_BURSTWRAP_H           (85),
		.PKT_BURSTWRAP_L           (80),
		.PKT_BYTE_CNT_H            (79),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (106),
		.PKT_PROTECTION_L          (104),
		.PKT_RESPONSE_STATUS_H     (112),
		.PKT_RESPONSE_STATUS_L     (111),
		.PKT_BURST_SIZE_H          (88),
		.PKT_BURST_SIZE_L          (86),
		.ST_CHANNEL_W              (12),
		.ST_DATA_W                 (113),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                  //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                           //       clk_reset.reset
		.m0_address              (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_009_src_ready),                                                               //              cp.ready
		.cp_valid                (cmd_xbar_mux_009_src_valid),                                                               //                .valid
		.cp_data                 (cmd_xbar_mux_009_src_data),                                                                //                .data
		.cp_startofpacket        (cmd_xbar_mux_009_src_startofpacket),                                                       //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_009_src_endofpacket),                                                         //                .endofpacket
		.cp_channel              (cmd_xbar_mux_009_src_channel),                                                             //                .channel
		.rf_sink_ready           (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (114),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                  //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                           // clk_reset.reset
		.in_data           (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                    // (terminated)
		.csr_read          (1'b0),                                                                                     // (terminated)
		.csr_write         (1'b0),                                                                                     // (terminated)
		.csr_readdata      (),                                                                                         // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                     // (terminated)
		.almost_full_data  (),                                                                                         // (terminated)
		.almost_empty_data (),                                                                                         // (terminated)
		.in_empty          (1'b0),                                                                                     // (terminated)
		.out_empty         (),                                                                                         // (terminated)
		.in_error          (1'b0),                                                                                     // (terminated)
		.out_error         (),                                                                                         // (terminated)
		.in_channel        (1'b0),                                                                                     // (terminated)
		.out_channel       ()                                                                                          // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (93),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (98),
		.PKT_SRC_ID_L              (95),
		.PKT_DEST_ID_H             (102),
		.PKT_DEST_ID_L             (99),
		.PKT_BURSTWRAP_H           (85),
		.PKT_BURSTWRAP_L           (80),
		.PKT_BYTE_CNT_H            (79),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (106),
		.PKT_PROTECTION_L          (104),
		.PKT_RESPONSE_STATUS_H     (112),
		.PKT_RESPONSE_STATUS_L     (111),
		.PKT_BURST_SIZE_H          (88),
		.PKT_BURST_SIZE_L          (86),
		.ST_CHANNEL_W              (12),
		.ST_DATA_W                 (113),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) jtaguart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                           //             clk.clk
		.reset                   (rst_controller_002_reset_out_reset),                                                                //       clk_reset.reset
		.m0_address              (jtaguart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (jtaguart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (jtaguart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (jtaguart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (jtaguart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (jtaguart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (jtaguart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (jtaguart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (jtaguart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (jtaguart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (jtaguart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (jtaguart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (jtaguart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (jtaguart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (jtaguart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (jtaguart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_002_src3_ready),                                                                     //              cp.ready
		.cp_valid                (cmd_xbar_demux_002_src3_valid),                                                                     //                .valid
		.cp_data                 (cmd_xbar_demux_002_src3_data),                                                                      //                .data
		.cp_startofpacket        (cmd_xbar_demux_002_src3_startofpacket),                                                             //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_002_src3_endofpacket),                                                               //                .endofpacket
		.cp_channel              (cmd_xbar_demux_002_src3_channel),                                                                   //                .channel
		.rf_sink_ready           (jtaguart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (jtaguart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (jtaguart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (jtaguart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (jtaguart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (jtaguart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (jtaguart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (jtaguart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (jtaguart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (jtaguart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (jtaguart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (jtaguart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (jtaguart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (jtaguart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (jtaguart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (jtaguart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (114),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) jtaguart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                           //       clk.clk
		.reset             (rst_controller_002_reset_out_reset),                                                                // clk_reset.reset
		.in_data           (jtaguart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (jtaguart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (jtaguart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (jtaguart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (jtaguart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (jtaguart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (jtaguart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (jtaguart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (jtaguart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (jtaguart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                             // (terminated)
		.csr_read          (1'b0),                                                                                              // (terminated)
		.csr_write         (1'b0),                                                                                              // (terminated)
		.csr_readdata      (),                                                                                                  // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                              // (terminated)
		.almost_full_data  (),                                                                                                  // (terminated)
		.almost_empty_data (),                                                                                                  // (terminated)
		.in_empty          (1'b0),                                                                                              // (terminated)
		.out_empty         (),                                                                                                  // (terminated)
		.in_error          (1'b0),                                                                                              // (terminated)
		.out_error         (),                                                                                                  // (terminated)
		.in_channel        (1'b0),                                                                                              // (terminated)
		.out_channel       ()                                                                                                   // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (93),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (98),
		.PKT_SRC_ID_L              (95),
		.PKT_DEST_ID_H             (102),
		.PKT_DEST_ID_L             (99),
		.PKT_BURSTWRAP_H           (85),
		.PKT_BURSTWRAP_L           (80),
		.PKT_BYTE_CNT_H            (79),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (106),
		.PKT_PROTECTION_L          (104),
		.PKT_RESPONSE_STATUS_H     (112),
		.PKT_RESPONSE_STATUS_L     (111),
		.PKT_BURST_SIZE_H          (88),
		.PKT_BURST_SIZE_L          (86),
		.ST_CHANNEL_W              (12),
		.ST_DATA_W                 (113),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) prio_arbiter_0_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                         //       clk_reset.reset
		.m0_address              (prio_arbiter_0_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (prio_arbiter_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (prio_arbiter_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (prio_arbiter_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (prio_arbiter_0_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (prio_arbiter_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (prio_arbiter_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (prio_arbiter_0_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (prio_arbiter_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (prio_arbiter_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (prio_arbiter_0_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (prio_arbiter_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (prio_arbiter_0_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (prio_arbiter_0_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (prio_arbiter_0_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (prio_arbiter_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_002_src4_ready),                                                          //              cp.ready
		.cp_valid                (cmd_xbar_demux_002_src4_valid),                                                          //                .valid
		.cp_data                 (cmd_xbar_demux_002_src4_data),                                                           //                .data
		.cp_startofpacket        (cmd_xbar_demux_002_src4_startofpacket),                                                  //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_002_src4_endofpacket),                                                    //                .endofpacket
		.cp_channel              (cmd_xbar_demux_002_src4_channel),                                                        //                .channel
		.rf_sink_ready           (prio_arbiter_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (prio_arbiter_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (prio_arbiter_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (prio_arbiter_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (prio_arbiter_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (prio_arbiter_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (prio_arbiter_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (prio_arbiter_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (prio_arbiter_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (prio_arbiter_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (prio_arbiter_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (prio_arbiter_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (prio_arbiter_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (prio_arbiter_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (prio_arbiter_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (prio_arbiter_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (114),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) prio_arbiter_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                         // clk_reset.reset
		.in_data           (prio_arbiter_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (prio_arbiter_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (prio_arbiter_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (prio_arbiter_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (prio_arbiter_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (prio_arbiter_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (prio_arbiter_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (prio_arbiter_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (prio_arbiter_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (prio_arbiter_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                  // (terminated)
		.csr_read          (1'b0),                                                                                   // (terminated)
		.csr_write         (1'b0),                                                                                   // (terminated)
		.csr_readdata      (),                                                                                       // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                   // (terminated)
		.almost_full_data  (),                                                                                       // (terminated)
		.almost_empty_data (),                                                                                       // (terminated)
		.in_empty          (1'b0),                                                                                   // (terminated)
		.out_empty         (),                                                                                       // (terminated)
		.in_error          (1'b0),                                                                                   // (terminated)
		.out_error         (),                                                                                       // (terminated)
		.in_channel        (1'b0),                                                                                   // (terminated)
		.out_channel       ()                                                                                        // (terminated)
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (96),
		.PKT_PROTECTION_L          (94),
		.PKT_BEGIN_BURST           (89),
		.PKT_BURSTWRAP_H           (81),
		.PKT_BURSTWRAP_L           (76),
		.PKT_BURST_SIZE_H          (84),
		.PKT_BURST_SIZE_L          (82),
		.PKT_BURST_TYPE_H          (86),
		.PKT_BURST_TYPE_L          (85),
		.PKT_BYTE_CNT_H            (75),
		.PKT_BYTE_CNT_L            (70),
		.PKT_ADDR_H                (63),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (64),
		.PKT_TRANS_POSTED          (65),
		.PKT_TRANS_WRITE           (66),
		.PKT_TRANS_READ            (67),
		.PKT_TRANS_LOCK            (68),
		.PKT_TRANS_EXCLUSIVE       (69),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (91),
		.PKT_SRC_ID_L              (91),
		.PKT_DEST_ID_H             (92),
		.PKT_DEST_ID_L             (92),
		.PKT_THREAD_ID_H           (93),
		.PKT_THREAD_ID_L           (93),
		.PKT_CACHE_H               (100),
		.PKT_CACHE_L               (97),
		.PKT_DATA_SIDEBAND_H       (88),
		.PKT_DATA_SIDEBAND_L       (88),
		.PKT_QOS_H                 (90),
		.PKT_QOS_L                 (90),
		.PKT_ADDR_SIDEBAND_H       (87),
		.PKT_ADDR_SIDEBAND_L       (87),
		.ST_DATA_W                 (103),
		.ST_CHANNEL_W              (1),
		.AV_BURSTCOUNT_W           (6),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (0),
		.BURSTWRAP_VALUE           (63),
		.CACHE_VALUE               (4'b0000)
	) traffic_gen_0_avalon_master_0_translator_avalon_universal_master_0_agent (
		.clk              (clk_clk),                                                                                   //       clk.clk
		.reset            (rst_controller_reset_out_reset),                                                            // clk_reset.reset
		.av_address       (traffic_gen_0_avalon_master_0_translator_avalon_universal_master_0_address),                //        av.address
		.av_write         (traffic_gen_0_avalon_master_0_translator_avalon_universal_master_0_write),                  //          .write
		.av_read          (traffic_gen_0_avalon_master_0_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata     (traffic_gen_0_avalon_master_0_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata      (traffic_gen_0_avalon_master_0_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest   (traffic_gen_0_avalon_master_0_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid (traffic_gen_0_avalon_master_0_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable    (traffic_gen_0_avalon_master_0_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount    (traffic_gen_0_avalon_master_0_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess   (traffic_gen_0_avalon_master_0_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock          (traffic_gen_0_avalon_master_0_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid         (traffic_gen_0_avalon_master_0_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data          (traffic_gen_0_avalon_master_0_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket (traffic_gen_0_avalon_master_0_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket   (traffic_gen_0_avalon_master_0_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready         (traffic_gen_0_avalon_master_0_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid         (rsp_xbar_demux_012_src0_valid),                                                             //        rp.valid
		.rp_data          (rsp_xbar_demux_012_src0_data),                                                              //          .data
		.rp_channel       (rsp_xbar_demux_012_src0_channel),                                                           //          .channel
		.rp_startofpacket (rsp_xbar_demux_012_src0_startofpacket),                                                     //          .startofpacket
		.rp_endofpacket   (rsp_xbar_demux_012_src0_endofpacket),                                                       //          .endofpacket
		.rp_ready         (rsp_xbar_demux_012_src0_ready)                                                              //          .ready
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (89),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (63),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (64),
		.PKT_TRANS_POSTED          (65),
		.PKT_TRANS_WRITE           (66),
		.PKT_TRANS_READ            (67),
		.PKT_TRANS_LOCK            (68),
		.PKT_SRC_ID_H              (91),
		.PKT_SRC_ID_L              (91),
		.PKT_DEST_ID_H             (92),
		.PKT_DEST_ID_L             (92),
		.PKT_BURSTWRAP_H           (81),
		.PKT_BURSTWRAP_L           (76),
		.PKT_BYTE_CNT_H            (75),
		.PKT_BYTE_CNT_L            (70),
		.PKT_PROTECTION_H          (96),
		.PKT_PROTECTION_L          (94),
		.PKT_RESPONSE_STATUS_H     (102),
		.PKT_RESPONSE_STATUS_L     (101),
		.PKT_BURST_SIZE_H          (84),
		.PKT_BURST_SIZE_L          (82),
		.ST_CHANNEL_W              (1),
		.ST_DATA_W                 (103),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) prio_arbiter_0_s2_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                         //       clk_reset.reset
		.m0_address              (prio_arbiter_0_s2_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (prio_arbiter_0_s2_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (prio_arbiter_0_s2_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (prio_arbiter_0_s2_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (prio_arbiter_0_s2_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (prio_arbiter_0_s2_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (prio_arbiter_0_s2_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (prio_arbiter_0_s2_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (prio_arbiter_0_s2_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (prio_arbiter_0_s2_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (prio_arbiter_0_s2_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (prio_arbiter_0_s2_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (prio_arbiter_0_s2_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (prio_arbiter_0_s2_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (prio_arbiter_0_s2_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (prio_arbiter_0_s2_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (burst_adapter_008_source0_ready),                                                        //              cp.ready
		.cp_valid                (burst_adapter_008_source0_valid),                                                        //                .valid
		.cp_data                 (burst_adapter_008_source0_data),                                                         //                .data
		.cp_startofpacket        (burst_adapter_008_source0_startofpacket),                                                //                .startofpacket
		.cp_endofpacket          (burst_adapter_008_source0_endofpacket),                                                  //                .endofpacket
		.cp_channel              (burst_adapter_008_source0_channel),                                                      //                .channel
		.rf_sink_ready           (prio_arbiter_0_s2_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (prio_arbiter_0_s2_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (prio_arbiter_0_s2_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (prio_arbiter_0_s2_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (prio_arbiter_0_s2_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (prio_arbiter_0_s2_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (prio_arbiter_0_s2_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (prio_arbiter_0_s2_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (prio_arbiter_0_s2_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (prio_arbiter_0_s2_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (prio_arbiter_0_s2_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (prio_arbiter_0_s2_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (prio_arbiter_0_s2_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (prio_arbiter_0_s2_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (prio_arbiter_0_s2_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (prio_arbiter_0_s2_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (104),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) prio_arbiter_0_s2_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                         // clk_reset.reset
		.in_data           (prio_arbiter_0_s2_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (prio_arbiter_0_s2_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (prio_arbiter_0_s2_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (prio_arbiter_0_s2_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (prio_arbiter_0_s2_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (prio_arbiter_0_s2_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (prio_arbiter_0_s2_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (prio_arbiter_0_s2_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (prio_arbiter_0_s2_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (prio_arbiter_0_s2_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                  // (terminated)
		.csr_read          (1'b0),                                                                                   // (terminated)
		.csr_write         (1'b0),                                                                                   // (terminated)
		.csr_readdata      (),                                                                                       // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                   // (terminated)
		.almost_full_data  (),                                                                                       // (terminated)
		.almost_empty_data (),                                                                                       // (terminated)
		.in_empty          (1'b0),                                                                                   // (terminated)
		.out_empty         (),                                                                                       // (terminated)
		.in_error          (1'b0),                                                                                   // (terminated)
		.out_error         (),                                                                                       // (terminated)
		.in_channel        (1'b0),                                                                                   // (terminated)
		.out_channel       ()                                                                                        // (terminated)
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (96),
		.PKT_PROTECTION_L          (94),
		.PKT_BEGIN_BURST           (89),
		.PKT_BURSTWRAP_H           (81),
		.PKT_BURSTWRAP_L           (76),
		.PKT_BURST_SIZE_H          (84),
		.PKT_BURST_SIZE_L          (82),
		.PKT_BURST_TYPE_H          (86),
		.PKT_BURST_TYPE_L          (85),
		.PKT_BYTE_CNT_H            (75),
		.PKT_BYTE_CNT_L            (70),
		.PKT_ADDR_H                (63),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (64),
		.PKT_TRANS_POSTED          (65),
		.PKT_TRANS_WRITE           (66),
		.PKT_TRANS_READ            (67),
		.PKT_TRANS_LOCK            (68),
		.PKT_TRANS_EXCLUSIVE       (69),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (91),
		.PKT_SRC_ID_L              (91),
		.PKT_DEST_ID_H             (92),
		.PKT_DEST_ID_L             (92),
		.PKT_THREAD_ID_H           (93),
		.PKT_THREAD_ID_L           (93),
		.PKT_CACHE_H               (100),
		.PKT_CACHE_L               (97),
		.PKT_DATA_SIDEBAND_H       (88),
		.PKT_DATA_SIDEBAND_L       (88),
		.PKT_QOS_H                 (90),
		.PKT_QOS_L                 (90),
		.PKT_ADDR_SIDEBAND_H       (87),
		.PKT_ADDR_SIDEBAND_L       (87),
		.ST_DATA_W                 (103),
		.ST_CHANNEL_W              (1),
		.AV_BURSTCOUNT_W           (6),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (0),
		.BURSTWRAP_VALUE           (63),
		.CACHE_VALUE               (4'b0000)
	) traffic_gen_1_avalon_master_0_translator_avalon_universal_master_0_agent (
		.clk              (clk_clk),                                                                                   //       clk.clk
		.reset            (rst_controller_reset_out_reset),                                                            // clk_reset.reset
		.av_address       (traffic_gen_1_avalon_master_0_translator_avalon_universal_master_0_address),                //        av.address
		.av_write         (traffic_gen_1_avalon_master_0_translator_avalon_universal_master_0_write),                  //          .write
		.av_read          (traffic_gen_1_avalon_master_0_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata     (traffic_gen_1_avalon_master_0_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata      (traffic_gen_1_avalon_master_0_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest   (traffic_gen_1_avalon_master_0_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid (traffic_gen_1_avalon_master_0_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable    (traffic_gen_1_avalon_master_0_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount    (traffic_gen_1_avalon_master_0_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess   (traffic_gen_1_avalon_master_0_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock          (traffic_gen_1_avalon_master_0_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid         (traffic_gen_1_avalon_master_0_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data          (traffic_gen_1_avalon_master_0_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket (traffic_gen_1_avalon_master_0_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket   (traffic_gen_1_avalon_master_0_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready         (traffic_gen_1_avalon_master_0_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid         (rsp_xbar_demux_013_src0_valid),                                                             //        rp.valid
		.rp_data          (rsp_xbar_demux_013_src0_data),                                                              //          .data
		.rp_channel       (rsp_xbar_demux_013_src0_channel),                                                           //          .channel
		.rp_startofpacket (rsp_xbar_demux_013_src0_startofpacket),                                                     //          .startofpacket
		.rp_endofpacket   (rsp_xbar_demux_013_src0_endofpacket),                                                       //          .endofpacket
		.rp_ready         (rsp_xbar_demux_013_src0_ready)                                                              //          .ready
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (89),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (63),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (64),
		.PKT_TRANS_POSTED          (65),
		.PKT_TRANS_WRITE           (66),
		.PKT_TRANS_READ            (67),
		.PKT_TRANS_LOCK            (68),
		.PKT_SRC_ID_H              (91),
		.PKT_SRC_ID_L              (91),
		.PKT_DEST_ID_H             (92),
		.PKT_DEST_ID_L             (92),
		.PKT_BURSTWRAP_H           (81),
		.PKT_BURSTWRAP_L           (76),
		.PKT_BYTE_CNT_H            (75),
		.PKT_BYTE_CNT_L            (70),
		.PKT_PROTECTION_H          (96),
		.PKT_PROTECTION_L          (94),
		.PKT_RESPONSE_STATUS_H     (102),
		.PKT_RESPONSE_STATUS_L     (101),
		.PKT_BURST_SIZE_H          (84),
		.PKT_BURST_SIZE_L          (82),
		.ST_CHANNEL_W              (1),
		.ST_DATA_W                 (103),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) prio_arbiter_0_s3_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                         //       clk_reset.reset
		.m0_address              (prio_arbiter_0_s3_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (prio_arbiter_0_s3_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (prio_arbiter_0_s3_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (prio_arbiter_0_s3_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (prio_arbiter_0_s3_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (prio_arbiter_0_s3_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (prio_arbiter_0_s3_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (prio_arbiter_0_s3_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (prio_arbiter_0_s3_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (prio_arbiter_0_s3_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (prio_arbiter_0_s3_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (prio_arbiter_0_s3_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (prio_arbiter_0_s3_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (prio_arbiter_0_s3_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (prio_arbiter_0_s3_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (prio_arbiter_0_s3_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (burst_adapter_009_source0_ready),                                                        //              cp.ready
		.cp_valid                (burst_adapter_009_source0_valid),                                                        //                .valid
		.cp_data                 (burst_adapter_009_source0_data),                                                         //                .data
		.cp_startofpacket        (burst_adapter_009_source0_startofpacket),                                                //                .startofpacket
		.cp_endofpacket          (burst_adapter_009_source0_endofpacket),                                                  //                .endofpacket
		.cp_channel              (burst_adapter_009_source0_channel),                                                      //                .channel
		.rf_sink_ready           (prio_arbiter_0_s3_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (prio_arbiter_0_s3_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (prio_arbiter_0_s3_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (prio_arbiter_0_s3_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (prio_arbiter_0_s3_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (prio_arbiter_0_s3_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (prio_arbiter_0_s3_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (prio_arbiter_0_s3_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (prio_arbiter_0_s3_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (prio_arbiter_0_s3_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (prio_arbiter_0_s3_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (prio_arbiter_0_s3_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (prio_arbiter_0_s3_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (prio_arbiter_0_s3_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (prio_arbiter_0_s3_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (prio_arbiter_0_s3_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (104),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) prio_arbiter_0_s3_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                         // clk_reset.reset
		.in_data           (prio_arbiter_0_s3_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (prio_arbiter_0_s3_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (prio_arbiter_0_s3_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (prio_arbiter_0_s3_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (prio_arbiter_0_s3_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (prio_arbiter_0_s3_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (prio_arbiter_0_s3_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (prio_arbiter_0_s3_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (prio_arbiter_0_s3_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (prio_arbiter_0_s3_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                  // (terminated)
		.csr_read          (1'b0),                                                                                   // (terminated)
		.csr_write         (1'b0),                                                                                   // (terminated)
		.csr_readdata      (),                                                                                       // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                   // (terminated)
		.almost_full_data  (),                                                                                       // (terminated)
		.almost_empty_data (),                                                                                       // (terminated)
		.in_empty          (1'b0),                                                                                   // (terminated)
		.out_empty         (),                                                                                       // (terminated)
		.in_error          (1'b0),                                                                                   // (terminated)
		.out_error         (),                                                                                       // (terminated)
		.in_channel        (1'b0),                                                                                   // (terminated)
		.out_channel       ()                                                                                        // (terminated)
	);

	nios_system_addr_router addr_router (
		.sink_ready         (com_nios_instruction_master_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (com_nios_instruction_master_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (com_nios_instruction_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (com_nios_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (com_nios_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                                 //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                          // clk_reset.reset
		.src_ready          (addr_router_src_ready),                                                                   //       src.ready
		.src_valid          (addr_router_src_valid),                                                                   //          .valid
		.src_data           (addr_router_src_data),                                                                    //          .data
		.src_channel        (addr_router_src_channel),                                                                 //          .channel
		.src_startofpacket  (addr_router_src_startofpacket),                                                           //          .startofpacket
		.src_endofpacket    (addr_router_src_endofpacket)                                                              //          .endofpacket
	);

	nios_system_addr_router_001 addr_router_001 (
		.sink_ready         (com_nios_data_master_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (com_nios_data_master_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (com_nios_data_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (com_nios_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (com_nios_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                          //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                   // clk_reset.reset
		.src_ready          (addr_router_001_src_ready),                                                        //       src.ready
		.src_valid          (addr_router_001_src_valid),                                                        //          .valid
		.src_data           (addr_router_001_src_data),                                                         //          .data
		.src_channel        (addr_router_001_src_channel),                                                      //          .channel
		.src_startofpacket  (addr_router_001_src_startofpacket),                                                //          .startofpacket
		.src_endofpacket    (addr_router_001_src_endofpacket)                                                   //          .endofpacket
	);

	nios_system_addr_router_002 addr_router_002 (
		.sink_ready         (carcontrol_nios_data_master_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (carcontrol_nios_data_master_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (carcontrol_nios_data_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (carcontrol_nios_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (carcontrol_nios_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                                 //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                          // clk_reset.reset
		.src_ready          (addr_router_002_src_ready),                                                               //       src.ready
		.src_valid          (addr_router_002_src_valid),                                                               //          .valid
		.src_data           (addr_router_002_src_data),                                                                //          .data
		.src_channel        (addr_router_002_src_channel),                                                             //          .channel
		.src_startofpacket  (addr_router_002_src_startofpacket),                                                       //          .startofpacket
		.src_endofpacket    (addr_router_002_src_endofpacket)                                                          //          .endofpacket
	);

	nios_system_addr_router_003 addr_router_003 (
		.sink_ready         (carcontrol_nios_instruction_master_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (carcontrol_nios_instruction_master_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (carcontrol_nios_instruction_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (carcontrol_nios_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (carcontrol_nios_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                                        //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                                 // clk_reset.reset
		.src_ready          (addr_router_003_src_ready),                                                                      //       src.ready
		.src_valid          (addr_router_003_src_valid),                                                                      //          .valid
		.src_data           (addr_router_003_src_data),                                                                       //          .data
		.src_channel        (addr_router_003_src_channel),                                                                    //          .channel
		.src_startofpacket  (addr_router_003_src_startofpacket),                                                              //          .startofpacket
		.src_endofpacket    (addr_router_003_src_endofpacket)                                                                 //          .endofpacket
	);

	nios_system_addr_router_004 addr_router_004 (
		.sink_ready         (ethernet_subsystem_sgdma_rx_m_write_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (ethernet_subsystem_sgdma_rx_m_write_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (ethernet_subsystem_sgdma_rx_m_write_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (ethernet_subsystem_sgdma_rx_m_write_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (ethernet_subsystem_sgdma_rx_m_write_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                                         //       clk.clk
		.reset              (rst_controller_002_reset_out_reset),                                                              // clk_reset.reset
		.src_ready          (addr_router_004_src_ready),                                                                       //       src.ready
		.src_valid          (addr_router_004_src_valid),                                                                       //          .valid
		.src_data           (addr_router_004_src_data),                                                                        //          .data
		.src_channel        (addr_router_004_src_channel),                                                                     //          .channel
		.src_startofpacket  (addr_router_004_src_startofpacket),                                                               //          .startofpacket
		.src_endofpacket    (addr_router_004_src_endofpacket)                                                                  //          .endofpacket
	);

	nios_system_addr_router_004 addr_router_005 (
		.sink_ready         (ethernet_subsystem_sgdma_tx_m_read_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (ethernet_subsystem_sgdma_tx_m_read_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (ethernet_subsystem_sgdma_tx_m_read_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (ethernet_subsystem_sgdma_tx_m_read_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (ethernet_subsystem_sgdma_tx_m_read_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                                        //       clk.clk
		.reset              (rst_controller_002_reset_out_reset),                                                             // clk_reset.reset
		.src_ready          (addr_router_005_src_ready),                                                                      //       src.ready
		.src_valid          (addr_router_005_src_valid),                                                                      //          .valid
		.src_data           (addr_router_005_src_data),                                                                       //          .data
		.src_channel        (addr_router_005_src_channel),                                                                    //          .channel
		.src_startofpacket  (addr_router_005_src_startofpacket),                                                              //          .startofpacket
		.src_endofpacket    (addr_router_005_src_endofpacket)                                                                 //          .endofpacket
	);

	nios_system_id_router id_router (
		.sink_ready         (com_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (com_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (com_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (com_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (com_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                        // clk_reset.reset
		.src_ready          (id_router_src_ready),                                                                   //       src.ready
		.src_valid          (id_router_src_valid),                                                                   //          .valid
		.src_data           (id_router_src_data),                                                                    //          .data
		.src_channel        (id_router_src_channel),                                                                 //          .channel
		.src_startofpacket  (id_router_src_startofpacket),                                                           //          .startofpacket
		.src_endofpacket    (id_router_src_endofpacket)                                                              //          .endofpacket
	);

	nios_system_id_router_001 id_router_001 (
		.sink_ready         (com_memory_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (com_memory_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (com_memory_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (com_memory_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (com_memory_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                  //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                           // clk_reset.reset
		.src_ready          (id_router_001_src_ready),                                                  //       src.ready
		.src_valid          (id_router_001_src_valid),                                                  //          .valid
		.src_data           (id_router_001_src_data),                                                   //          .data
		.src_channel        (id_router_001_src_channel),                                                //          .channel
		.src_startofpacket  (id_router_001_src_startofpacket),                                          //          .startofpacket
		.src_endofpacket    (id_router_001_src_endofpacket)                                             //          .endofpacket
	);

	nios_system_id_router_002 id_router_002 (
		.sink_ready         (jtaguart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (jtaguart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (jtaguart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (jtaguart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (jtaguart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                                 //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                                      // clk_reset.reset
		.src_ready          (id_router_002_src_ready),                                                                 //       src.ready
		.src_valid          (id_router_002_src_valid),                                                                 //          .valid
		.src_data           (id_router_002_src_data),                                                                  //          .data
		.src_channel        (id_router_002_src_channel),                                                               //          .channel
		.src_startofpacket  (id_router_002_src_startofpacket),                                                         //          .startofpacket
		.src_endofpacket    (id_router_002_src_endofpacket)                                                            //          .endofpacket
	);

	nios_system_id_router_003 id_router_003 (
		.sink_ready         (shared_memory_mutex_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (shared_memory_mutex_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (shared_memory_mutex_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (shared_memory_mutex_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (shared_memory_mutex_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                           //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                    // clk_reset.reset
		.src_ready          (id_router_003_src_ready),                                                           //       src.ready
		.src_valid          (id_router_003_src_valid),                                                           //          .valid
		.src_data           (id_router_003_src_data),                                                            //          .data
		.src_channel        (id_router_003_src_channel),                                                         //          .channel
		.src_startofpacket  (id_router_003_src_startofpacket),                                                   //          .startofpacket
		.src_endofpacket    (id_router_003_src_endofpacket)                                                      //          .endofpacket
	);

	nios_system_id_router_002 id_router_004 (
		.sink_ready         (com_timer_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (com_timer_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (com_timer_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (com_timer_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (com_timer_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                 //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                          // clk_reset.reset
		.src_ready          (id_router_004_src_ready),                                                 //       src.ready
		.src_valid          (id_router_004_src_valid),                                                 //          .valid
		.src_data           (id_router_004_src_data),                                                  //          .data
		.src_channel        (id_router_004_src_channel),                                               //          .channel
		.src_startofpacket  (id_router_004_src_startofpacket),                                         //          .startofpacket
		.src_endofpacket    (id_router_004_src_endofpacket)                                            //          .endofpacket
	);

	nios_system_id_router_002 id_router_005 (
		.sink_ready         (ethernet_subsystem_ethernet_bridge_s0_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (ethernet_subsystem_ethernet_bridge_s0_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (ethernet_subsystem_ethernet_bridge_s0_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (ethernet_subsystem_ethernet_bridge_s0_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (ethernet_subsystem_ethernet_bridge_s0_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                                          //       clk.clk
		.reset              (rst_controller_002_reset_out_reset),                                                               // clk_reset.reset
		.src_ready          (id_router_005_src_ready),                                                                          //       src.ready
		.src_valid          (id_router_005_src_valid),                                                                          //          .valid
		.src_data           (id_router_005_src_data),                                                                           //          .data
		.src_channel        (id_router_005_src_channel),                                                                        //          .channel
		.src_startofpacket  (id_router_005_src_startofpacket),                                                                  //          .startofpacket
		.src_endofpacket    (id_router_005_src_endofpacket)                                                                     //          .endofpacket
	);

	nios_system_id_router_002 id_router_006 (
		.sink_ready         (ethernet_subsystem_descriptor_memory_s2_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (ethernet_subsystem_descriptor_memory_s2_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (ethernet_subsystem_descriptor_memory_s2_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (ethernet_subsystem_descriptor_memory_s2_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (ethernet_subsystem_descriptor_memory_s2_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                                            //       clk.clk
		.reset              (rst_controller_002_reset_out_reset),                                                                 // clk_reset.reset
		.src_ready          (id_router_006_src_ready),                                                                            //       src.ready
		.src_valid          (id_router_006_src_valid),                                                                            //          .valid
		.src_data           (id_router_006_src_data),                                                                             //          .data
		.src_channel        (id_router_006_src_channel),                                                                          //          .channel
		.src_startofpacket  (id_router_006_src_startofpacket),                                                                    //          .startofpacket
		.src_endofpacket    (id_router_006_src_endofpacket)                                                                       //          .endofpacket
	);

	nios_system_id_router_002 id_router_007 (
		.sink_ready         (prio_arbiter_0_s0_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (prio_arbiter_0_s0_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (prio_arbiter_0_s0_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (prio_arbiter_0_s0_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (prio_arbiter_0_s0_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                      //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                               // clk_reset.reset
		.src_ready          (id_router_007_src_ready),                                                      //       src.ready
		.src_valid          (id_router_007_src_valid),                                                      //          .valid
		.src_data           (id_router_007_src_data),                                                       //          .data
		.src_channel        (id_router_007_src_channel),                                                    //          .channel
		.src_startofpacket  (id_router_007_src_startofpacket),                                              //          .startofpacket
		.src_endofpacket    (id_router_007_src_endofpacket)                                                 //          .endofpacket
	);

	nios_system_id_router_008 id_router_008 (
		.sink_ready         (carcontrol_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (carcontrol_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (carcontrol_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (carcontrol_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (carcontrol_nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                                      //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                               // clk_reset.reset
		.src_ready          (id_router_008_src_ready),                                                                      //       src.ready
		.src_valid          (id_router_008_src_valid),                                                                      //          .valid
		.src_data           (id_router_008_src_data),                                                                       //          .data
		.src_channel        (id_router_008_src_channel),                                                                    //          .channel
		.src_startofpacket  (id_router_008_src_startofpacket),                                                              //          .startofpacket
		.src_endofpacket    (id_router_008_src_endofpacket)                                                                 //          .endofpacket
	);

	nios_system_id_router_008 id_router_009 (
		.sink_ready         (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                        //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                 // clk_reset.reset
		.src_ready          (id_router_009_src_ready),                                                        //       src.ready
		.src_valid          (id_router_009_src_valid),                                                        //          .valid
		.src_data           (id_router_009_src_data),                                                         //          .data
		.src_channel        (id_router_009_src_channel),                                                      //          .channel
		.src_startofpacket  (id_router_009_src_startofpacket),                                                //          .startofpacket
		.src_endofpacket    (id_router_009_src_endofpacket)                                                   //          .endofpacket
	);

	nios_system_id_router_010 id_router_010 (
		.sink_ready         (jtaguart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (jtaguart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (jtaguart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (jtaguart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (jtaguart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                                 //       clk.clk
		.reset              (rst_controller_002_reset_out_reset),                                                      // clk_reset.reset
		.src_ready          (id_router_010_src_ready),                                                                 //       src.ready
		.src_valid          (id_router_010_src_valid),                                                                 //          .valid
		.src_data           (id_router_010_src_data),                                                                  //          .data
		.src_channel        (id_router_010_src_channel),                                                               //          .channel
		.src_startofpacket  (id_router_010_src_startofpacket),                                                         //          .startofpacket
		.src_endofpacket    (id_router_010_src_endofpacket)                                                            //          .endofpacket
	);

	nios_system_id_router_010 id_router_011 (
		.sink_ready         (prio_arbiter_0_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (prio_arbiter_0_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (prio_arbiter_0_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (prio_arbiter_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (prio_arbiter_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                      //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                               // clk_reset.reset
		.src_ready          (id_router_011_src_ready),                                                      //       src.ready
		.src_valid          (id_router_011_src_valid),                                                      //          .valid
		.src_data           (id_router_011_src_data),                                                       //          .data
		.src_channel        (id_router_011_src_channel),                                                    //          .channel
		.src_startofpacket  (id_router_011_src_startofpacket),                                              //          .startofpacket
		.src_endofpacket    (id_router_011_src_endofpacket)                                                 //          .endofpacket
	);

	nios_system_addr_router_006 addr_router_006 (
		.sink_ready         (traffic_gen_0_avalon_master_0_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (traffic_gen_0_avalon_master_0_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (traffic_gen_0_avalon_master_0_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (traffic_gen_0_avalon_master_0_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (traffic_gen_0_avalon_master_0_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                                   //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                            // clk_reset.reset
		.src_ready          (addr_router_006_src_ready),                                                                 //       src.ready
		.src_valid          (addr_router_006_src_valid),                                                                 //          .valid
		.src_data           (addr_router_006_src_data),                                                                  //          .data
		.src_channel        (addr_router_006_src_channel),                                                               //          .channel
		.src_startofpacket  (addr_router_006_src_startofpacket),                                                         //          .startofpacket
		.src_endofpacket    (addr_router_006_src_endofpacket)                                                            //          .endofpacket
	);

	nios_system_id_router_012 id_router_012 (
		.sink_ready         (prio_arbiter_0_s2_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (prio_arbiter_0_s2_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (prio_arbiter_0_s2_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (prio_arbiter_0_s2_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (prio_arbiter_0_s2_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                      //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                               // clk_reset.reset
		.src_ready          (id_router_012_src_ready),                                                      //       src.ready
		.src_valid          (id_router_012_src_valid),                                                      //          .valid
		.src_data           (id_router_012_src_data),                                                       //          .data
		.src_channel        (id_router_012_src_channel),                                                    //          .channel
		.src_startofpacket  (id_router_012_src_startofpacket),                                              //          .startofpacket
		.src_endofpacket    (id_router_012_src_endofpacket)                                                 //          .endofpacket
	);

	nios_system_addr_router_006 addr_router_007 (
		.sink_ready         (traffic_gen_1_avalon_master_0_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (traffic_gen_1_avalon_master_0_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (traffic_gen_1_avalon_master_0_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (traffic_gen_1_avalon_master_0_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (traffic_gen_1_avalon_master_0_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                                   //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                            // clk_reset.reset
		.src_ready          (addr_router_007_src_ready),                                                                 //       src.ready
		.src_valid          (addr_router_007_src_valid),                                                                 //          .valid
		.src_data           (addr_router_007_src_data),                                                                  //          .data
		.src_channel        (addr_router_007_src_channel),                                                               //          .channel
		.src_startofpacket  (addr_router_007_src_startofpacket),                                                         //          .startofpacket
		.src_endofpacket    (addr_router_007_src_endofpacket)                                                            //          .endofpacket
	);

	nios_system_id_router_012 id_router_013 (
		.sink_ready         (prio_arbiter_0_s3_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (prio_arbiter_0_s3_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (prio_arbiter_0_s3_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (prio_arbiter_0_s3_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (prio_arbiter_0_s3_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                      //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                               // clk_reset.reset
		.src_ready          (id_router_013_src_ready),                                                      //       src.ready
		.src_valid          (id_router_013_src_valid),                                                      //          .valid
		.src_data           (id_router_013_src_data),                                                       //          .data
		.src_channel        (id_router_013_src_channel),                                                    //          .channel
		.src_startofpacket  (id_router_013_src_startofpacket),                                              //          .startofpacket
		.src_endofpacket    (id_router_013_src_endofpacket)                                                 //          .endofpacket
	);

	altera_merlin_traffic_limiter #(
		.PKT_DEST_ID_H             (102),
		.PKT_DEST_ID_L             (99),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.MAX_OUTSTANDING_RESPONSES (9),
		.PIPELINED                 (0),
		.ST_DATA_W                 (113),
		.ST_CHANNEL_W              (12),
		.VALID_WIDTH               (12),
		.ENFORCE_ORDER             (1),
		.PREVENT_HAZARDS           (0),
		.PKT_BYTE_CNT_H            (79),
		.PKT_BYTE_CNT_L            (74),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32)
	) limiter (
		.clk                    (clk_clk),                        //       clk.clk
		.reset                  (rst_controller_reset_out_reset), // clk_reset.reset
		.cmd_sink_ready         (addr_router_src_ready),          //  cmd_sink.ready
		.cmd_sink_valid         (addr_router_src_valid),          //          .valid
		.cmd_sink_data          (addr_router_src_data),           //          .data
		.cmd_sink_channel       (addr_router_src_channel),        //          .channel
		.cmd_sink_startofpacket (addr_router_src_startofpacket),  //          .startofpacket
		.cmd_sink_endofpacket   (addr_router_src_endofpacket),    //          .endofpacket
		.cmd_src_ready          (limiter_cmd_src_ready),          //   cmd_src.ready
		.cmd_src_data           (limiter_cmd_src_data),           //          .data
		.cmd_src_channel        (limiter_cmd_src_channel),        //          .channel
		.cmd_src_startofpacket  (limiter_cmd_src_startofpacket),  //          .startofpacket
		.cmd_src_endofpacket    (limiter_cmd_src_endofpacket),    //          .endofpacket
		.rsp_sink_ready         (rsp_xbar_mux_src_ready),         //  rsp_sink.ready
		.rsp_sink_valid         (rsp_xbar_mux_src_valid),         //          .valid
		.rsp_sink_channel       (rsp_xbar_mux_src_channel),       //          .channel
		.rsp_sink_data          (rsp_xbar_mux_src_data),          //          .data
		.rsp_sink_startofpacket (rsp_xbar_mux_src_startofpacket), //          .startofpacket
		.rsp_sink_endofpacket   (rsp_xbar_mux_src_endofpacket),   //          .endofpacket
		.rsp_src_ready          (limiter_rsp_src_ready),          //   rsp_src.ready
		.rsp_src_valid          (limiter_rsp_src_valid),          //          .valid
		.rsp_src_data           (limiter_rsp_src_data),           //          .data
		.rsp_src_channel        (limiter_rsp_src_channel),        //          .channel
		.rsp_src_startofpacket  (limiter_rsp_src_startofpacket),  //          .startofpacket
		.rsp_src_endofpacket    (limiter_rsp_src_endofpacket),    //          .endofpacket
		.cmd_src_valid          (limiter_cmd_valid_data)          // cmd_valid.data
	);

	altera_merlin_traffic_limiter #(
		.PKT_DEST_ID_H             (102),
		.PKT_DEST_ID_L             (99),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.MAX_OUTSTANDING_RESPONSES (9),
		.PIPELINED                 (0),
		.ST_DATA_W                 (113),
		.ST_CHANNEL_W              (12),
		.VALID_WIDTH               (12),
		.ENFORCE_ORDER             (1),
		.PREVENT_HAZARDS           (0),
		.PKT_BYTE_CNT_H            (79),
		.PKT_BYTE_CNT_L            (74),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32)
	) limiter_001 (
		.clk                    (clk_clk),                            //       clk.clk
		.reset                  (rst_controller_reset_out_reset),     // clk_reset.reset
		.cmd_sink_ready         (addr_router_001_src_ready),          //  cmd_sink.ready
		.cmd_sink_valid         (addr_router_001_src_valid),          //          .valid
		.cmd_sink_data          (addr_router_001_src_data),           //          .data
		.cmd_sink_channel       (addr_router_001_src_channel),        //          .channel
		.cmd_sink_startofpacket (addr_router_001_src_startofpacket),  //          .startofpacket
		.cmd_sink_endofpacket   (addr_router_001_src_endofpacket),    //          .endofpacket
		.cmd_src_ready          (limiter_001_cmd_src_ready),          //   cmd_src.ready
		.cmd_src_data           (limiter_001_cmd_src_data),           //          .data
		.cmd_src_channel        (limiter_001_cmd_src_channel),        //          .channel
		.cmd_src_startofpacket  (limiter_001_cmd_src_startofpacket),  //          .startofpacket
		.cmd_src_endofpacket    (limiter_001_cmd_src_endofpacket),    //          .endofpacket
		.rsp_sink_ready         (rsp_xbar_mux_001_src_ready),         //  rsp_sink.ready
		.rsp_sink_valid         (rsp_xbar_mux_001_src_valid),         //          .valid
		.rsp_sink_channel       (rsp_xbar_mux_001_src_channel),       //          .channel
		.rsp_sink_data          (rsp_xbar_mux_001_src_data),          //          .data
		.rsp_sink_startofpacket (rsp_xbar_mux_001_src_startofpacket), //          .startofpacket
		.rsp_sink_endofpacket   (rsp_xbar_mux_001_src_endofpacket),   //          .endofpacket
		.rsp_src_ready          (limiter_001_rsp_src_ready),          //   rsp_src.ready
		.rsp_src_valid          (limiter_001_rsp_src_valid),          //          .valid
		.rsp_src_data           (limiter_001_rsp_src_data),           //          .data
		.rsp_src_channel        (limiter_001_rsp_src_channel),        //          .channel
		.rsp_src_startofpacket  (limiter_001_rsp_src_startofpacket),  //          .startofpacket
		.rsp_src_endofpacket    (limiter_001_rsp_src_endofpacket),    //          .endofpacket
		.cmd_src_valid          (limiter_001_cmd_valid_data)          // cmd_valid.data
	);

	altera_merlin_traffic_limiter #(
		.PKT_DEST_ID_H             (102),
		.PKT_DEST_ID_L             (99),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.MAX_OUTSTANDING_RESPONSES (1),
		.PIPELINED                 (0),
		.ST_DATA_W                 (113),
		.ST_CHANNEL_W              (12),
		.VALID_WIDTH               (12),
		.ENFORCE_ORDER             (1),
		.PREVENT_HAZARDS           (0),
		.PKT_BYTE_CNT_H            (79),
		.PKT_BYTE_CNT_L            (74),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32)
	) limiter_002 (
		.clk                    (clk_clk),                            //       clk.clk
		.reset                  (rst_controller_reset_out_reset),     // clk_reset.reset
		.cmd_sink_ready         (addr_router_003_src_ready),          //  cmd_sink.ready
		.cmd_sink_valid         (addr_router_003_src_valid),          //          .valid
		.cmd_sink_data          (addr_router_003_src_data),           //          .data
		.cmd_sink_channel       (addr_router_003_src_channel),        //          .channel
		.cmd_sink_startofpacket (addr_router_003_src_startofpacket),  //          .startofpacket
		.cmd_sink_endofpacket   (addr_router_003_src_endofpacket),    //          .endofpacket
		.cmd_src_ready          (limiter_002_cmd_src_ready),          //   cmd_src.ready
		.cmd_src_data           (limiter_002_cmd_src_data),           //          .data
		.cmd_src_channel        (limiter_002_cmd_src_channel),        //          .channel
		.cmd_src_startofpacket  (limiter_002_cmd_src_startofpacket),  //          .startofpacket
		.cmd_src_endofpacket    (limiter_002_cmd_src_endofpacket),    //          .endofpacket
		.rsp_sink_ready         (rsp_xbar_mux_003_src_ready),         //  rsp_sink.ready
		.rsp_sink_valid         (rsp_xbar_mux_003_src_valid),         //          .valid
		.rsp_sink_channel       (rsp_xbar_mux_003_src_channel),       //          .channel
		.rsp_sink_data          (rsp_xbar_mux_003_src_data),          //          .data
		.rsp_sink_startofpacket (rsp_xbar_mux_003_src_startofpacket), //          .startofpacket
		.rsp_sink_endofpacket   (rsp_xbar_mux_003_src_endofpacket),   //          .endofpacket
		.rsp_src_ready          (limiter_002_rsp_src_ready),          //   rsp_src.ready
		.rsp_src_valid          (limiter_002_rsp_src_valid),          //          .valid
		.rsp_src_data           (limiter_002_rsp_src_data),           //          .data
		.rsp_src_channel        (limiter_002_rsp_src_channel),        //          .channel
		.rsp_src_startofpacket  (limiter_002_rsp_src_startofpacket),  //          .startofpacket
		.rsp_src_endofpacket    (limiter_002_rsp_src_endofpacket),    //          .endofpacket
		.cmd_src_valid          (limiter_002_cmd_valid_data)          // cmd_valid.data
	);

	altera_merlin_burst_adapter #(
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_BEGIN_BURST           (93),
		.PKT_BYTE_CNT_H            (79),
		.PKT_BYTE_CNT_L            (74),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_BURST_SIZE_H          (88),
		.PKT_BURST_SIZE_L          (86),
		.PKT_BURST_TYPE_H          (90),
		.PKT_BURST_TYPE_L          (89),
		.PKT_BURSTWRAP_H           (85),
		.PKT_BURSTWRAP_L           (80),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.OUT_NARROW_SIZE           (0),
		.IN_NARROW_SIZE            (0),
		.OUT_FIXED                 (0),
		.OUT_COMPLETE_WRAP         (0),
		.ST_DATA_W                 (113),
		.ST_CHANNEL_W              (12),
		.OUT_BYTE_CNT_H            (76),
		.OUT_BURSTWRAP_H           (85),
		.COMPRESSED_READ_SUPPORT   (1),
		.BYTEENABLE_SYNTHESIS      (0),
		.PIPE_INPUTS               (0),
		.NO_WRAP_SUPPORT           (0),
		.BURSTWRAP_CONST_MASK      (31),
		.BURSTWRAP_CONST_VALUE     (31)
	) burst_adapter (
		.clk                   (clk_clk),                             //       cr0.clk
		.reset                 (rst_controller_reset_out_reset),      // cr0_reset.reset
		.sink0_valid           (cmd_xbar_mux_src_valid),              //     sink0.valid
		.sink0_data            (cmd_xbar_mux_src_data),               //          .data
		.sink0_channel         (cmd_xbar_mux_src_channel),            //          .channel
		.sink0_startofpacket   (cmd_xbar_mux_src_startofpacket),      //          .startofpacket
		.sink0_endofpacket     (cmd_xbar_mux_src_endofpacket),        //          .endofpacket
		.sink0_ready           (cmd_xbar_mux_src_ready),              //          .ready
		.source0_valid         (burst_adapter_source0_valid),         //   source0.valid
		.source0_data          (burst_adapter_source0_data),          //          .data
		.source0_channel       (burst_adapter_source0_channel),       //          .channel
		.source0_startofpacket (burst_adapter_source0_startofpacket), //          .startofpacket
		.source0_endofpacket   (burst_adapter_source0_endofpacket),   //          .endofpacket
		.source0_ready         (burst_adapter_source0_ready)          //          .ready
	);

	altera_merlin_burst_adapter #(
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_BEGIN_BURST           (93),
		.PKT_BYTE_CNT_H            (79),
		.PKT_BYTE_CNT_L            (74),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_BURST_SIZE_H          (88),
		.PKT_BURST_SIZE_L          (86),
		.PKT_BURST_TYPE_H          (90),
		.PKT_BURST_TYPE_L          (89),
		.PKT_BURSTWRAP_H           (85),
		.PKT_BURSTWRAP_L           (80),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.OUT_NARROW_SIZE           (0),
		.IN_NARROW_SIZE            (0),
		.OUT_FIXED                 (0),
		.OUT_COMPLETE_WRAP         (0),
		.ST_DATA_W                 (113),
		.ST_CHANNEL_W              (12),
		.OUT_BYTE_CNT_H            (76),
		.OUT_BURSTWRAP_H           (85),
		.COMPRESSED_READ_SUPPORT   (1),
		.BYTEENABLE_SYNTHESIS      (0),
		.PIPE_INPUTS               (0),
		.NO_WRAP_SUPPORT           (0),
		.BURSTWRAP_CONST_MASK      (31),
		.BURSTWRAP_CONST_VALUE     (31)
	) burst_adapter_001 (
		.clk                   (clk_clk),                                 //       cr0.clk
		.reset                 (rst_controller_reset_out_reset),          // cr0_reset.reset
		.sink0_valid           (cmd_xbar_mux_001_src_valid),              //     sink0.valid
		.sink0_data            (cmd_xbar_mux_001_src_data),               //          .data
		.sink0_channel         (cmd_xbar_mux_001_src_channel),            //          .channel
		.sink0_startofpacket   (cmd_xbar_mux_001_src_startofpacket),      //          .startofpacket
		.sink0_endofpacket     (cmd_xbar_mux_001_src_endofpacket),        //          .endofpacket
		.sink0_ready           (cmd_xbar_mux_001_src_ready),              //          .ready
		.source0_valid         (burst_adapter_001_source0_valid),         //   source0.valid
		.source0_data          (burst_adapter_001_source0_data),          //          .data
		.source0_channel       (burst_adapter_001_source0_channel),       //          .channel
		.source0_startofpacket (burst_adapter_001_source0_startofpacket), //          .startofpacket
		.source0_endofpacket   (burst_adapter_001_source0_endofpacket),   //          .endofpacket
		.source0_ready         (burst_adapter_001_source0_ready)          //          .ready
	);

	altera_merlin_burst_adapter #(
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_BEGIN_BURST           (93),
		.PKT_BYTE_CNT_H            (79),
		.PKT_BYTE_CNT_L            (74),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_BURST_SIZE_H          (88),
		.PKT_BURST_SIZE_L          (86),
		.PKT_BURST_TYPE_H          (90),
		.PKT_BURST_TYPE_L          (89),
		.PKT_BURSTWRAP_H           (85),
		.PKT_BURSTWRAP_L           (80),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.OUT_NARROW_SIZE           (0),
		.IN_NARROW_SIZE            (0),
		.OUT_FIXED                 (0),
		.OUT_COMPLETE_WRAP         (0),
		.ST_DATA_W                 (113),
		.ST_CHANNEL_W              (12),
		.OUT_BYTE_CNT_H            (76),
		.OUT_BURSTWRAP_H           (85),
		.COMPRESSED_READ_SUPPORT   (1),
		.BYTEENABLE_SYNTHESIS      (0),
		.PIPE_INPUTS               (0),
		.NO_WRAP_SUPPORT           (0),
		.BURSTWRAP_CONST_MASK      (63),
		.BURSTWRAP_CONST_VALUE     (63)
	) burst_adapter_002 (
		.clk                   (clk_clk),                                 //       cr0.clk
		.reset                 (rst_controller_001_reset_out_reset),      // cr0_reset.reset
		.sink0_valid           (cmd_xbar_demux_001_src2_valid),           //     sink0.valid
		.sink0_data            (cmd_xbar_demux_001_src2_data),            //          .data
		.sink0_channel         (cmd_xbar_demux_001_src2_channel),         //          .channel
		.sink0_startofpacket   (cmd_xbar_demux_001_src2_startofpacket),   //          .startofpacket
		.sink0_endofpacket     (cmd_xbar_demux_001_src2_endofpacket),     //          .endofpacket
		.sink0_ready           (cmd_xbar_demux_001_src2_ready),           //          .ready
		.source0_valid         (burst_adapter_002_source0_valid),         //   source0.valid
		.source0_data          (burst_adapter_002_source0_data),          //          .data
		.source0_channel       (burst_adapter_002_source0_channel),       //          .channel
		.source0_startofpacket (burst_adapter_002_source0_startofpacket), //          .startofpacket
		.source0_endofpacket   (burst_adapter_002_source0_endofpacket),   //          .endofpacket
		.source0_ready         (burst_adapter_002_source0_ready)          //          .ready
	);

	altera_merlin_burst_adapter #(
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_BEGIN_BURST           (93),
		.PKT_BYTE_CNT_H            (79),
		.PKT_BYTE_CNT_L            (74),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_BURST_SIZE_H          (88),
		.PKT_BURST_SIZE_L          (86),
		.PKT_BURST_TYPE_H          (90),
		.PKT_BURST_TYPE_L          (89),
		.PKT_BURSTWRAP_H           (85),
		.PKT_BURSTWRAP_L           (80),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.OUT_NARROW_SIZE           (0),
		.IN_NARROW_SIZE            (0),
		.OUT_FIXED                 (0),
		.OUT_COMPLETE_WRAP         (0),
		.ST_DATA_W                 (113),
		.ST_CHANNEL_W              (12),
		.OUT_BYTE_CNT_H            (76),
		.OUT_BURSTWRAP_H           (85),
		.COMPRESSED_READ_SUPPORT   (1),
		.BYTEENABLE_SYNTHESIS      (0),
		.PIPE_INPUTS               (0),
		.NO_WRAP_SUPPORT           (0),
		.BURSTWRAP_CONST_MASK      (63),
		.BURSTWRAP_CONST_VALUE     (63)
	) burst_adapter_003 (
		.clk                   (clk_clk),                                 //       cr0.clk
		.reset                 (rst_controller_reset_out_reset),          // cr0_reset.reset
		.sink0_valid           (cmd_xbar_mux_003_src_valid),              //     sink0.valid
		.sink0_data            (cmd_xbar_mux_003_src_data),               //          .data
		.sink0_channel         (cmd_xbar_mux_003_src_channel),            //          .channel
		.sink0_startofpacket   (cmd_xbar_mux_003_src_startofpacket),      //          .startofpacket
		.sink0_endofpacket     (cmd_xbar_mux_003_src_endofpacket),        //          .endofpacket
		.sink0_ready           (cmd_xbar_mux_003_src_ready),              //          .ready
		.source0_valid         (burst_adapter_003_source0_valid),         //   source0.valid
		.source0_data          (burst_adapter_003_source0_data),          //          .data
		.source0_channel       (burst_adapter_003_source0_channel),       //          .channel
		.source0_startofpacket (burst_adapter_003_source0_startofpacket), //          .startofpacket
		.source0_endofpacket   (burst_adapter_003_source0_endofpacket),   //          .endofpacket
		.source0_ready         (burst_adapter_003_source0_ready)          //          .ready
	);

	altera_merlin_burst_adapter #(
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_BEGIN_BURST           (93),
		.PKT_BYTE_CNT_H            (79),
		.PKT_BYTE_CNT_L            (74),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_BURST_SIZE_H          (88),
		.PKT_BURST_SIZE_L          (86),
		.PKT_BURST_TYPE_H          (90),
		.PKT_BURST_TYPE_L          (89),
		.PKT_BURSTWRAP_H           (85),
		.PKT_BURSTWRAP_L           (80),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.OUT_NARROW_SIZE           (0),
		.IN_NARROW_SIZE            (0),
		.OUT_FIXED                 (0),
		.OUT_COMPLETE_WRAP         (0),
		.ST_DATA_W                 (113),
		.ST_CHANNEL_W              (12),
		.OUT_BYTE_CNT_H            (76),
		.OUT_BURSTWRAP_H           (85),
		.COMPRESSED_READ_SUPPORT   (1),
		.BYTEENABLE_SYNTHESIS      (0),
		.PIPE_INPUTS               (0),
		.NO_WRAP_SUPPORT           (0),
		.BURSTWRAP_CONST_MASK      (63),
		.BURSTWRAP_CONST_VALUE     (63)
	) burst_adapter_004 (
		.clk                   (clk_clk),                                 //       cr0.clk
		.reset                 (rst_controller_reset_out_reset),          // cr0_reset.reset
		.sink0_valid           (cmd_xbar_demux_001_src4_valid),           //     sink0.valid
		.sink0_data            (cmd_xbar_demux_001_src4_data),            //          .data
		.sink0_channel         (cmd_xbar_demux_001_src4_channel),         //          .channel
		.sink0_startofpacket   (cmd_xbar_demux_001_src4_startofpacket),   //          .startofpacket
		.sink0_endofpacket     (cmd_xbar_demux_001_src4_endofpacket),     //          .endofpacket
		.sink0_ready           (cmd_xbar_demux_001_src4_ready),           //          .ready
		.source0_valid         (burst_adapter_004_source0_valid),         //   source0.valid
		.source0_data          (burst_adapter_004_source0_data),          //          .data
		.source0_channel       (burst_adapter_004_source0_channel),       //          .channel
		.source0_startofpacket (burst_adapter_004_source0_startofpacket), //          .startofpacket
		.source0_endofpacket   (burst_adapter_004_source0_endofpacket),   //          .endofpacket
		.source0_ready         (burst_adapter_004_source0_ready)          //          .ready
	);

	altera_merlin_burst_adapter #(
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_BEGIN_BURST           (93),
		.PKT_BYTE_CNT_H            (79),
		.PKT_BYTE_CNT_L            (74),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_BURST_SIZE_H          (88),
		.PKT_BURST_SIZE_L          (86),
		.PKT_BURST_TYPE_H          (90),
		.PKT_BURST_TYPE_L          (89),
		.PKT_BURSTWRAP_H           (85),
		.PKT_BURSTWRAP_L           (80),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.OUT_NARROW_SIZE           (0),
		.IN_NARROW_SIZE            (0),
		.OUT_FIXED                 (0),
		.OUT_COMPLETE_WRAP         (0),
		.ST_DATA_W                 (113),
		.ST_CHANNEL_W              (12),
		.OUT_BYTE_CNT_H            (76),
		.OUT_BURSTWRAP_H           (85),
		.COMPRESSED_READ_SUPPORT   (1),
		.BYTEENABLE_SYNTHESIS      (0),
		.PIPE_INPUTS               (0),
		.NO_WRAP_SUPPORT           (0),
		.BURSTWRAP_CONST_MASK      (63),
		.BURSTWRAP_CONST_VALUE     (63)
	) burst_adapter_005 (
		.clk                   (clk_clk),                                 //       cr0.clk
		.reset                 (rst_controller_002_reset_out_reset),      // cr0_reset.reset
		.sink0_valid           (cmd_xbar_demux_001_src5_valid),           //     sink0.valid
		.sink0_data            (cmd_xbar_demux_001_src5_data),            //          .data
		.sink0_channel         (cmd_xbar_demux_001_src5_channel),         //          .channel
		.sink0_startofpacket   (cmd_xbar_demux_001_src5_startofpacket),   //          .startofpacket
		.sink0_endofpacket     (cmd_xbar_demux_001_src5_endofpacket),     //          .endofpacket
		.sink0_ready           (cmd_xbar_demux_001_src5_ready),           //          .ready
		.source0_valid         (burst_adapter_005_source0_valid),         //   source0.valid
		.source0_data          (burst_adapter_005_source0_data),          //          .data
		.source0_channel       (burst_adapter_005_source0_channel),       //          .channel
		.source0_startofpacket (burst_adapter_005_source0_startofpacket), //          .startofpacket
		.source0_endofpacket   (burst_adapter_005_source0_endofpacket),   //          .endofpacket
		.source0_ready         (burst_adapter_005_source0_ready)          //          .ready
	);

	altera_merlin_burst_adapter #(
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_BEGIN_BURST           (93),
		.PKT_BYTE_CNT_H            (79),
		.PKT_BYTE_CNT_L            (74),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_BURST_SIZE_H          (88),
		.PKT_BURST_SIZE_L          (86),
		.PKT_BURST_TYPE_H          (90),
		.PKT_BURST_TYPE_L          (89),
		.PKT_BURSTWRAP_H           (85),
		.PKT_BURSTWRAP_L           (80),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.OUT_NARROW_SIZE           (0),
		.IN_NARROW_SIZE            (0),
		.OUT_FIXED                 (0),
		.OUT_COMPLETE_WRAP         (0),
		.ST_DATA_W                 (113),
		.ST_CHANNEL_W              (12),
		.OUT_BYTE_CNT_H            (76),
		.OUT_BURSTWRAP_H           (85),
		.COMPRESSED_READ_SUPPORT   (1),
		.BYTEENABLE_SYNTHESIS      (0),
		.PIPE_INPUTS               (0),
		.NO_WRAP_SUPPORT           (0),
		.BURSTWRAP_CONST_MASK      (63),
		.BURSTWRAP_CONST_VALUE     (63)
	) burst_adapter_006 (
		.clk                   (clk_clk),                                 //       cr0.clk
		.reset                 (rst_controller_002_reset_out_reset),      // cr0_reset.reset
		.sink0_valid           (cmd_xbar_demux_001_src6_valid),           //     sink0.valid
		.sink0_data            (cmd_xbar_demux_001_src6_data),            //          .data
		.sink0_channel         (cmd_xbar_demux_001_src6_channel),         //          .channel
		.sink0_startofpacket   (cmd_xbar_demux_001_src6_startofpacket),   //          .startofpacket
		.sink0_endofpacket     (cmd_xbar_demux_001_src6_endofpacket),     //          .endofpacket
		.sink0_ready           (cmd_xbar_demux_001_src6_ready),           //          .ready
		.source0_valid         (burst_adapter_006_source0_valid),         //   source0.valid
		.source0_data          (burst_adapter_006_source0_data),          //          .data
		.source0_channel       (burst_adapter_006_source0_channel),       //          .channel
		.source0_startofpacket (burst_adapter_006_source0_startofpacket), //          .startofpacket
		.source0_endofpacket   (burst_adapter_006_source0_endofpacket),   //          .endofpacket
		.source0_ready         (burst_adapter_006_source0_ready)          //          .ready
	);

	altera_merlin_burst_adapter #(
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_BEGIN_BURST           (93),
		.PKT_BYTE_CNT_H            (79),
		.PKT_BYTE_CNT_L            (74),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_BURST_SIZE_H          (88),
		.PKT_BURST_SIZE_L          (86),
		.PKT_BURST_TYPE_H          (90),
		.PKT_BURST_TYPE_L          (89),
		.PKT_BURSTWRAP_H           (85),
		.PKT_BURSTWRAP_L           (80),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.OUT_NARROW_SIZE           (0),
		.IN_NARROW_SIZE            (0),
		.OUT_FIXED                 (0),
		.OUT_COMPLETE_WRAP         (0),
		.ST_DATA_W                 (113),
		.ST_CHANNEL_W              (12),
		.OUT_BYTE_CNT_H            (76),
		.OUT_BURSTWRAP_H           (85),
		.COMPRESSED_READ_SUPPORT   (1),
		.BYTEENABLE_SYNTHESIS      (0),
		.PIPE_INPUTS               (0),
		.NO_WRAP_SUPPORT           (0),
		.BURSTWRAP_CONST_MASK      (63),
		.BURSTWRAP_CONST_VALUE     (63)
	) burst_adapter_007 (
		.clk                   (clk_clk),                                 //       cr0.clk
		.reset                 (rst_controller_reset_out_reset),          // cr0_reset.reset
		.sink0_valid           (cmd_xbar_demux_001_src7_valid),           //     sink0.valid
		.sink0_data            (cmd_xbar_demux_001_src7_data),            //          .data
		.sink0_channel         (cmd_xbar_demux_001_src7_channel),         //          .channel
		.sink0_startofpacket   (cmd_xbar_demux_001_src7_startofpacket),   //          .startofpacket
		.sink0_endofpacket     (cmd_xbar_demux_001_src7_endofpacket),     //          .endofpacket
		.sink0_ready           (cmd_xbar_demux_001_src7_ready),           //          .ready
		.source0_valid         (burst_adapter_007_source0_valid),         //   source0.valid
		.source0_data          (burst_adapter_007_source0_data),          //          .data
		.source0_channel       (burst_adapter_007_source0_channel),       //          .channel
		.source0_startofpacket (burst_adapter_007_source0_startofpacket), //          .startofpacket
		.source0_endofpacket   (burst_adapter_007_source0_endofpacket),   //          .endofpacket
		.source0_ready         (burst_adapter_007_source0_ready)          //          .ready
	);

	altera_merlin_burst_adapter #(
		.PKT_ADDR_H                (63),
		.PKT_ADDR_L                (36),
		.PKT_BEGIN_BURST           (89),
		.PKT_BYTE_CNT_H            (75),
		.PKT_BYTE_CNT_L            (70),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_BURST_SIZE_H          (84),
		.PKT_BURST_SIZE_L          (82),
		.PKT_BURST_TYPE_H          (86),
		.PKT_BURST_TYPE_L          (85),
		.PKT_BURSTWRAP_H           (81),
		.PKT_BURSTWRAP_L           (76),
		.PKT_TRANS_COMPRESSED_READ (64),
		.PKT_TRANS_WRITE           (66),
		.PKT_TRANS_READ            (67),
		.OUT_NARROW_SIZE           (0),
		.IN_NARROW_SIZE            (0),
		.OUT_FIXED                 (0),
		.OUT_COMPLETE_WRAP         (0),
		.ST_DATA_W                 (103),
		.ST_CHANNEL_W              (1),
		.OUT_BYTE_CNT_H            (72),
		.OUT_BURSTWRAP_H           (81),
		.COMPRESSED_READ_SUPPORT   (1),
		.BYTEENABLE_SYNTHESIS      (0),
		.PIPE_INPUTS               (0),
		.NO_WRAP_SUPPORT           (0),
		.BURSTWRAP_CONST_MASK      (63),
		.BURSTWRAP_CONST_VALUE     (63)
	) burst_adapter_008 (
		.clk                   (clk_clk),                                 //       cr0.clk
		.reset                 (rst_controller_reset_out_reset),          // cr0_reset.reset
		.sink0_valid           (cmd_xbar_demux_006_src0_valid),           //     sink0.valid
		.sink0_data            (cmd_xbar_demux_006_src0_data),            //          .data
		.sink0_channel         (cmd_xbar_demux_006_src0_channel),         //          .channel
		.sink0_startofpacket   (cmd_xbar_demux_006_src0_startofpacket),   //          .startofpacket
		.sink0_endofpacket     (cmd_xbar_demux_006_src0_endofpacket),     //          .endofpacket
		.sink0_ready           (cmd_xbar_demux_006_src0_ready),           //          .ready
		.source0_valid         (burst_adapter_008_source0_valid),         //   source0.valid
		.source0_data          (burst_adapter_008_source0_data),          //          .data
		.source0_channel       (burst_adapter_008_source0_channel),       //          .channel
		.source0_startofpacket (burst_adapter_008_source0_startofpacket), //          .startofpacket
		.source0_endofpacket   (burst_adapter_008_source0_endofpacket),   //          .endofpacket
		.source0_ready         (burst_adapter_008_source0_ready)          //          .ready
	);

	altera_merlin_burst_adapter #(
		.PKT_ADDR_H                (63),
		.PKT_ADDR_L                (36),
		.PKT_BEGIN_BURST           (89),
		.PKT_BYTE_CNT_H            (75),
		.PKT_BYTE_CNT_L            (70),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_BURST_SIZE_H          (84),
		.PKT_BURST_SIZE_L          (82),
		.PKT_BURST_TYPE_H          (86),
		.PKT_BURST_TYPE_L          (85),
		.PKT_BURSTWRAP_H           (81),
		.PKT_BURSTWRAP_L           (76),
		.PKT_TRANS_COMPRESSED_READ (64),
		.PKT_TRANS_WRITE           (66),
		.PKT_TRANS_READ            (67),
		.OUT_NARROW_SIZE           (0),
		.IN_NARROW_SIZE            (0),
		.OUT_FIXED                 (0),
		.OUT_COMPLETE_WRAP         (0),
		.ST_DATA_W                 (103),
		.ST_CHANNEL_W              (1),
		.OUT_BYTE_CNT_H            (72),
		.OUT_BURSTWRAP_H           (81),
		.COMPRESSED_READ_SUPPORT   (1),
		.BYTEENABLE_SYNTHESIS      (0),
		.PIPE_INPUTS               (0),
		.NO_WRAP_SUPPORT           (0),
		.BURSTWRAP_CONST_MASK      (63),
		.BURSTWRAP_CONST_VALUE     (63)
	) burst_adapter_009 (
		.clk                   (clk_clk),                                 //       cr0.clk
		.reset                 (rst_controller_reset_out_reset),          // cr0_reset.reset
		.sink0_valid           (cmd_xbar_demux_007_src0_valid),           //     sink0.valid
		.sink0_data            (cmd_xbar_demux_007_src0_data),            //          .data
		.sink0_channel         (cmd_xbar_demux_007_src0_channel),         //          .channel
		.sink0_startofpacket   (cmd_xbar_demux_007_src0_startofpacket),   //          .startofpacket
		.sink0_endofpacket     (cmd_xbar_demux_007_src0_endofpacket),     //          .endofpacket
		.sink0_ready           (cmd_xbar_demux_007_src0_ready),           //          .ready
		.source0_valid         (burst_adapter_009_source0_valid),         //   source0.valid
		.source0_data          (burst_adapter_009_source0_data),          //          .data
		.source0_channel       (burst_adapter_009_source0_channel),       //          .channel
		.source0_startofpacket (burst_adapter_009_source0_startofpacket), //          .startofpacket
		.source0_endofpacket   (burst_adapter_009_source0_endofpacket),   //          .endofpacket
		.source0_ready         (burst_adapter_009_source0_ready)          //          .ready
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (3),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2)
	) rst_controller (
		.reset_in0  (~reset_reset_n),                                // reset_in0.reset
		.reset_in1  (com_nios_jtag_debug_module_reset_reset),        // reset_in1.reset
		.reset_in2  (carcontrol_nios_jtag_debug_module_reset_reset), // reset_in2.reset
		.clk        (clk_clk),                                       //       clk.clk
		.reset_out  (rst_controller_reset_out_reset),                // reset_out.reset
		.reset_in3  (1'b0),                                          // (terminated)
		.reset_in4  (1'b0),                                          // (terminated)
		.reset_in5  (1'b0),                                          // (terminated)
		.reset_in6  (1'b0),                                          // (terminated)
		.reset_in7  (1'b0),                                          // (terminated)
		.reset_in8  (1'b0),                                          // (terminated)
		.reset_in9  (1'b0),                                          // (terminated)
		.reset_in10 (1'b0),                                          // (terminated)
		.reset_in11 (1'b0),                                          // (terminated)
		.reset_in12 (1'b0),                                          // (terminated)
		.reset_in13 (1'b0),                                          // (terminated)
		.reset_in14 (1'b0),                                          // (terminated)
		.reset_in15 (1'b0)                                           // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (2),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2)
	) rst_controller_001 (
		.reset_in0  (~reset_reset_n),                         // reset_in0.reset
		.reset_in1  (com_nios_jtag_debug_module_reset_reset), // reset_in1.reset
		.clk        (clk_clk),                                //       clk.clk
		.reset_out  (rst_controller_001_reset_out_reset),     // reset_out.reset
		.reset_in2  (1'b0),                                   // (terminated)
		.reset_in3  (1'b0),                                   // (terminated)
		.reset_in4  (1'b0),                                   // (terminated)
		.reset_in5  (1'b0),                                   // (terminated)
		.reset_in6  (1'b0),                                   // (terminated)
		.reset_in7  (1'b0),                                   // (terminated)
		.reset_in8  (1'b0),                                   // (terminated)
		.reset_in9  (1'b0),                                   // (terminated)
		.reset_in10 (1'b0),                                   // (terminated)
		.reset_in11 (1'b0),                                   // (terminated)
		.reset_in12 (1'b0),                                   // (terminated)
		.reset_in13 (1'b0),                                   // (terminated)
		.reset_in14 (1'b0),                                   // (terminated)
		.reset_in15 (1'b0)                                    // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (1),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2)
	) rst_controller_002 (
		.reset_in0  (~reset_reset_n),                     // reset_in0.reset
		.clk        (clk_clk),                            //       clk.clk
		.reset_out  (rst_controller_002_reset_out_reset), // reset_out.reset
		.reset_in1  (1'b0),                               // (terminated)
		.reset_in2  (1'b0),                               // (terminated)
		.reset_in3  (1'b0),                               // (terminated)
		.reset_in4  (1'b0),                               // (terminated)
		.reset_in5  (1'b0),                               // (terminated)
		.reset_in6  (1'b0),                               // (terminated)
		.reset_in7  (1'b0),                               // (terminated)
		.reset_in8  (1'b0),                               // (terminated)
		.reset_in9  (1'b0),                               // (terminated)
		.reset_in10 (1'b0),                               // (terminated)
		.reset_in11 (1'b0),                               // (terminated)
		.reset_in12 (1'b0),                               // (terminated)
		.reset_in13 (1'b0),                               // (terminated)
		.reset_in14 (1'b0),                               // (terminated)
		.reset_in15 (1'b0)                                // (terminated)
	);

	nios_system_cmd_xbar_demux cmd_xbar_demux (
		.clk                (clk_clk),                           //        clk.clk
		.reset              (rst_controller_reset_out_reset),    //  clk_reset.reset
		.sink_ready         (limiter_cmd_src_ready),             //       sink.ready
		.sink_channel       (limiter_cmd_src_channel),           //           .channel
		.sink_data          (limiter_cmd_src_data),              //           .data
		.sink_startofpacket (limiter_cmd_src_startofpacket),     //           .startofpacket
		.sink_endofpacket   (limiter_cmd_src_endofpacket),       //           .endofpacket
		.sink_valid         (limiter_cmd_valid_data),            // sink_valid.data
		.src0_ready         (cmd_xbar_demux_src0_ready),         //       src0.ready
		.src0_valid         (cmd_xbar_demux_src0_valid),         //           .valid
		.src0_data          (cmd_xbar_demux_src0_data),          //           .data
		.src0_channel       (cmd_xbar_demux_src0_channel),       //           .channel
		.src0_startofpacket (cmd_xbar_demux_src0_startofpacket), //           .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_src0_endofpacket),   //           .endofpacket
		.src1_ready         (cmd_xbar_demux_src1_ready),         //       src1.ready
		.src1_valid         (cmd_xbar_demux_src1_valid),         //           .valid
		.src1_data          (cmd_xbar_demux_src1_data),          //           .data
		.src1_channel       (cmd_xbar_demux_src1_channel),       //           .channel
		.src1_startofpacket (cmd_xbar_demux_src1_startofpacket), //           .startofpacket
		.src1_endofpacket   (cmd_xbar_demux_src1_endofpacket)    //           .endofpacket
	);

	nios_system_cmd_xbar_demux_001 cmd_xbar_demux_001 (
		.clk                (clk_clk),                               //        clk.clk
		.reset              (rst_controller_reset_out_reset),        //  clk_reset.reset
		.sink_ready         (limiter_001_cmd_src_ready),             //       sink.ready
		.sink_channel       (limiter_001_cmd_src_channel),           //           .channel
		.sink_data          (limiter_001_cmd_src_data),              //           .data
		.sink_startofpacket (limiter_001_cmd_src_startofpacket),     //           .startofpacket
		.sink_endofpacket   (limiter_001_cmd_src_endofpacket),       //           .endofpacket
		.sink_valid         (limiter_001_cmd_valid_data),            // sink_valid.data
		.src0_ready         (cmd_xbar_demux_001_src0_ready),         //       src0.ready
		.src0_valid         (cmd_xbar_demux_001_src0_valid),         //           .valid
		.src0_data          (cmd_xbar_demux_001_src0_data),          //           .data
		.src0_channel       (cmd_xbar_demux_001_src0_channel),       //           .channel
		.src0_startofpacket (cmd_xbar_demux_001_src0_startofpacket), //           .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_001_src0_endofpacket),   //           .endofpacket
		.src1_ready         (cmd_xbar_demux_001_src1_ready),         //       src1.ready
		.src1_valid         (cmd_xbar_demux_001_src1_valid),         //           .valid
		.src1_data          (cmd_xbar_demux_001_src1_data),          //           .data
		.src1_channel       (cmd_xbar_demux_001_src1_channel),       //           .channel
		.src1_startofpacket (cmd_xbar_demux_001_src1_startofpacket), //           .startofpacket
		.src1_endofpacket   (cmd_xbar_demux_001_src1_endofpacket),   //           .endofpacket
		.src2_ready         (cmd_xbar_demux_001_src2_ready),         //       src2.ready
		.src2_valid         (cmd_xbar_demux_001_src2_valid),         //           .valid
		.src2_data          (cmd_xbar_demux_001_src2_data),          //           .data
		.src2_channel       (cmd_xbar_demux_001_src2_channel),       //           .channel
		.src2_startofpacket (cmd_xbar_demux_001_src2_startofpacket), //           .startofpacket
		.src2_endofpacket   (cmd_xbar_demux_001_src2_endofpacket),   //           .endofpacket
		.src3_ready         (cmd_xbar_demux_001_src3_ready),         //       src3.ready
		.src3_valid         (cmd_xbar_demux_001_src3_valid),         //           .valid
		.src3_data          (cmd_xbar_demux_001_src3_data),          //           .data
		.src3_channel       (cmd_xbar_demux_001_src3_channel),       //           .channel
		.src3_startofpacket (cmd_xbar_demux_001_src3_startofpacket), //           .startofpacket
		.src3_endofpacket   (cmd_xbar_demux_001_src3_endofpacket),   //           .endofpacket
		.src4_ready         (cmd_xbar_demux_001_src4_ready),         //       src4.ready
		.src4_valid         (cmd_xbar_demux_001_src4_valid),         //           .valid
		.src4_data          (cmd_xbar_demux_001_src4_data),          //           .data
		.src4_channel       (cmd_xbar_demux_001_src4_channel),       //           .channel
		.src4_startofpacket (cmd_xbar_demux_001_src4_startofpacket), //           .startofpacket
		.src4_endofpacket   (cmd_xbar_demux_001_src4_endofpacket),   //           .endofpacket
		.src5_ready         (cmd_xbar_demux_001_src5_ready),         //       src5.ready
		.src5_valid         (cmd_xbar_demux_001_src5_valid),         //           .valid
		.src5_data          (cmd_xbar_demux_001_src5_data),          //           .data
		.src5_channel       (cmd_xbar_demux_001_src5_channel),       //           .channel
		.src5_startofpacket (cmd_xbar_demux_001_src5_startofpacket), //           .startofpacket
		.src5_endofpacket   (cmd_xbar_demux_001_src5_endofpacket),   //           .endofpacket
		.src6_ready         (cmd_xbar_demux_001_src6_ready),         //       src6.ready
		.src6_valid         (cmd_xbar_demux_001_src6_valid),         //           .valid
		.src6_data          (cmd_xbar_demux_001_src6_data),          //           .data
		.src6_channel       (cmd_xbar_demux_001_src6_channel),       //           .channel
		.src6_startofpacket (cmd_xbar_demux_001_src6_startofpacket), //           .startofpacket
		.src6_endofpacket   (cmd_xbar_demux_001_src6_endofpacket),   //           .endofpacket
		.src7_ready         (cmd_xbar_demux_001_src7_ready),         //       src7.ready
		.src7_valid         (cmd_xbar_demux_001_src7_valid),         //           .valid
		.src7_data          (cmd_xbar_demux_001_src7_data),          //           .data
		.src7_channel       (cmd_xbar_demux_001_src7_channel),       //           .channel
		.src7_startofpacket (cmd_xbar_demux_001_src7_startofpacket), //           .startofpacket
		.src7_endofpacket   (cmd_xbar_demux_001_src7_endofpacket)    //           .endofpacket
	);

	nios_system_cmd_xbar_demux_002 cmd_xbar_demux_002 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (addr_router_002_src_ready),             //      sink.ready
		.sink_channel       (addr_router_002_src_channel),           //          .channel
		.sink_data          (addr_router_002_src_data),              //          .data
		.sink_startofpacket (addr_router_002_src_startofpacket),     //          .startofpacket
		.sink_endofpacket   (addr_router_002_src_endofpacket),       //          .endofpacket
		.sink_valid         (addr_router_002_src_valid),             //          .valid
		.src0_ready         (cmd_xbar_demux_002_src0_ready),         //      src0.ready
		.src0_valid         (cmd_xbar_demux_002_src0_valid),         //          .valid
		.src0_data          (cmd_xbar_demux_002_src0_data),          //          .data
		.src0_channel       (cmd_xbar_demux_002_src0_channel),       //          .channel
		.src0_startofpacket (cmd_xbar_demux_002_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_002_src0_endofpacket),   //          .endofpacket
		.src1_ready         (cmd_xbar_demux_002_src1_ready),         //      src1.ready
		.src1_valid         (cmd_xbar_demux_002_src1_valid),         //          .valid
		.src1_data          (cmd_xbar_demux_002_src1_data),          //          .data
		.src1_channel       (cmd_xbar_demux_002_src1_channel),       //          .channel
		.src1_startofpacket (cmd_xbar_demux_002_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (cmd_xbar_demux_002_src1_endofpacket),   //          .endofpacket
		.src2_ready         (cmd_xbar_demux_002_src2_ready),         //      src2.ready
		.src2_valid         (cmd_xbar_demux_002_src2_valid),         //          .valid
		.src2_data          (cmd_xbar_demux_002_src2_data),          //          .data
		.src2_channel       (cmd_xbar_demux_002_src2_channel),       //          .channel
		.src2_startofpacket (cmd_xbar_demux_002_src2_startofpacket), //          .startofpacket
		.src2_endofpacket   (cmd_xbar_demux_002_src2_endofpacket),   //          .endofpacket
		.src3_ready         (cmd_xbar_demux_002_src3_ready),         //      src3.ready
		.src3_valid         (cmd_xbar_demux_002_src3_valid),         //          .valid
		.src3_data          (cmd_xbar_demux_002_src3_data),          //          .data
		.src3_channel       (cmd_xbar_demux_002_src3_channel),       //          .channel
		.src3_startofpacket (cmd_xbar_demux_002_src3_startofpacket), //          .startofpacket
		.src3_endofpacket   (cmd_xbar_demux_002_src3_endofpacket),   //          .endofpacket
		.src4_ready         (cmd_xbar_demux_002_src4_ready),         //      src4.ready
		.src4_valid         (cmd_xbar_demux_002_src4_valid),         //          .valid
		.src4_data          (cmd_xbar_demux_002_src4_data),          //          .data
		.src4_channel       (cmd_xbar_demux_002_src4_channel),       //          .channel
		.src4_startofpacket (cmd_xbar_demux_002_src4_startofpacket), //          .startofpacket
		.src4_endofpacket   (cmd_xbar_demux_002_src4_endofpacket)    //          .endofpacket
	);

	nios_system_cmd_xbar_demux cmd_xbar_demux_003 (
		.clk                (clk_clk),                               //        clk.clk
		.reset              (rst_controller_reset_out_reset),        //  clk_reset.reset
		.sink_ready         (limiter_002_cmd_src_ready),             //       sink.ready
		.sink_channel       (limiter_002_cmd_src_channel),           //           .channel
		.sink_data          (limiter_002_cmd_src_data),              //           .data
		.sink_startofpacket (limiter_002_cmd_src_startofpacket),     //           .startofpacket
		.sink_endofpacket   (limiter_002_cmd_src_endofpacket),       //           .endofpacket
		.sink_valid         (limiter_002_cmd_valid_data),            // sink_valid.data
		.src0_ready         (cmd_xbar_demux_003_src0_ready),         //       src0.ready
		.src0_valid         (cmd_xbar_demux_003_src0_valid),         //           .valid
		.src0_data          (cmd_xbar_demux_003_src0_data),          //           .data
		.src0_channel       (cmd_xbar_demux_003_src0_channel),       //           .channel
		.src0_startofpacket (cmd_xbar_demux_003_src0_startofpacket), //           .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_003_src0_endofpacket),   //           .endofpacket
		.src1_ready         (cmd_xbar_demux_003_src1_ready),         //       src1.ready
		.src1_valid         (cmd_xbar_demux_003_src1_valid),         //           .valid
		.src1_data          (cmd_xbar_demux_003_src1_data),          //           .data
		.src1_channel       (cmd_xbar_demux_003_src1_channel),       //           .channel
		.src1_startofpacket (cmd_xbar_demux_003_src1_startofpacket), //           .startofpacket
		.src1_endofpacket   (cmd_xbar_demux_003_src1_endofpacket)    //           .endofpacket
	);

	nios_system_cmd_xbar_demux_004 cmd_xbar_demux_004 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_002_reset_out_reset),    // clk_reset.reset
		.sink_ready         (addr_router_004_src_ready),             //      sink.ready
		.sink_channel       (addr_router_004_src_channel),           //          .channel
		.sink_data          (addr_router_004_src_data),              //          .data
		.sink_startofpacket (addr_router_004_src_startofpacket),     //          .startofpacket
		.sink_endofpacket   (addr_router_004_src_endofpacket),       //          .endofpacket
		.sink_valid         (addr_router_004_src_valid),             //          .valid
		.src0_ready         (cmd_xbar_demux_004_src0_ready),         //      src0.ready
		.src0_valid         (cmd_xbar_demux_004_src0_valid),         //          .valid
		.src0_data          (cmd_xbar_demux_004_src0_data),          //          .data
		.src0_channel       (cmd_xbar_demux_004_src0_channel),       //          .channel
		.src0_startofpacket (cmd_xbar_demux_004_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_004_src0_endofpacket)    //          .endofpacket
	);

	nios_system_cmd_xbar_demux_004 cmd_xbar_demux_005 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_002_reset_out_reset),    // clk_reset.reset
		.sink_ready         (addr_router_005_src_ready),             //      sink.ready
		.sink_channel       (addr_router_005_src_channel),           //          .channel
		.sink_data          (addr_router_005_src_data),              //          .data
		.sink_startofpacket (addr_router_005_src_startofpacket),     //          .startofpacket
		.sink_endofpacket   (addr_router_005_src_endofpacket),       //          .endofpacket
		.sink_valid         (addr_router_005_src_valid),             //          .valid
		.src0_ready         (cmd_xbar_demux_005_src0_ready),         //      src0.ready
		.src0_valid         (cmd_xbar_demux_005_src0_valid),         //          .valid
		.src0_data          (cmd_xbar_demux_005_src0_data),          //          .data
		.src0_channel       (cmd_xbar_demux_005_src0_channel),       //          .channel
		.src0_startofpacket (cmd_xbar_demux_005_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_005_src0_endofpacket)    //          .endofpacket
	);

	nios_system_cmd_xbar_mux cmd_xbar_mux (
		.clk                 (clk_clk),                               //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (cmd_xbar_mux_src_ready),                //       src.ready
		.src_valid           (cmd_xbar_mux_src_valid),                //          .valid
		.src_data            (cmd_xbar_mux_src_data),                 //          .data
		.src_channel         (cmd_xbar_mux_src_channel),              //          .channel
		.src_startofpacket   (cmd_xbar_mux_src_startofpacket),        //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_src_endofpacket),          //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src0_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src0_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src0_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src0_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src0_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src0_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src0_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src0_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src0_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src0_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src0_endofpacket)    //          .endofpacket
	);

	nios_system_cmd_xbar_mux_001 cmd_xbar_mux_001 (
		.clk                 (clk_clk),                               //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (cmd_xbar_mux_001_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_001_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_001_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_001_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_001_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_001_src_endofpacket),      //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src1_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src1_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src1_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src1_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src1_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src1_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src1_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src1_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src1_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src1_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src1_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src1_endofpacket),   //          .endofpacket
		.sink2_ready         (cmd_xbar_demux_004_src0_ready),         //     sink2.ready
		.sink2_valid         (cmd_xbar_demux_004_src0_valid),         //          .valid
		.sink2_channel       (cmd_xbar_demux_004_src0_channel),       //          .channel
		.sink2_data          (cmd_xbar_demux_004_src0_data),          //          .data
		.sink2_startofpacket (cmd_xbar_demux_004_src0_startofpacket), //          .startofpacket
		.sink2_endofpacket   (cmd_xbar_demux_004_src0_endofpacket),   //          .endofpacket
		.sink3_ready         (cmd_xbar_demux_005_src0_ready),         //     sink3.ready
		.sink3_valid         (cmd_xbar_demux_005_src0_valid),         //          .valid
		.sink3_channel       (cmd_xbar_demux_005_src0_channel),       //          .channel
		.sink3_data          (cmd_xbar_demux_005_src0_data),          //          .data
		.sink3_startofpacket (cmd_xbar_demux_005_src0_startofpacket), //          .startofpacket
		.sink3_endofpacket   (cmd_xbar_demux_005_src0_endofpacket)    //          .endofpacket
	);

	nios_system_cmd_xbar_mux cmd_xbar_mux_003 (
		.clk                 (clk_clk),                               //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (cmd_xbar_mux_003_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_003_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_003_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_003_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_003_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_003_src_endofpacket),      //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_001_src3_ready),         //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_001_src3_valid),         //          .valid
		.sink0_channel       (cmd_xbar_demux_001_src3_channel),       //          .channel
		.sink0_data          (cmd_xbar_demux_001_src3_data),          //          .data
		.sink0_startofpacket (cmd_xbar_demux_001_src3_startofpacket), //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_001_src3_endofpacket),   //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_002_src0_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_002_src0_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_002_src0_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_002_src0_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_002_src0_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_002_src0_endofpacket)    //          .endofpacket
	);

	nios_system_cmd_xbar_mux cmd_xbar_mux_008 (
		.clk                 (clk_clk),                               //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (cmd_xbar_mux_008_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_008_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_008_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_008_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_008_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_008_src_endofpacket),      //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_002_src1_ready),         //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_002_src1_valid),         //          .valid
		.sink0_channel       (cmd_xbar_demux_002_src1_channel),       //          .channel
		.sink0_data          (cmd_xbar_demux_002_src1_data),          //          .data
		.sink0_startofpacket (cmd_xbar_demux_002_src1_startofpacket), //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_002_src1_endofpacket),   //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_003_src0_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_003_src0_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_003_src0_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_003_src0_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_003_src0_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_003_src0_endofpacket)    //          .endofpacket
	);

	nios_system_cmd_xbar_mux cmd_xbar_mux_009 (
		.clk                 (clk_clk),                               //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (cmd_xbar_mux_009_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_009_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_009_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_009_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_009_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_009_src_endofpacket),      //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_002_src2_ready),         //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_002_src2_valid),         //          .valid
		.sink0_channel       (cmd_xbar_demux_002_src2_channel),       //          .channel
		.sink0_data          (cmd_xbar_demux_002_src2_data),          //          .data
		.sink0_startofpacket (cmd_xbar_demux_002_src2_startofpacket), //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_002_src2_endofpacket),   //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_003_src1_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_003_src1_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_003_src1_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_003_src1_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_003_src1_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_003_src1_endofpacket)    //          .endofpacket
	);

	nios_system_rsp_xbar_demux rsp_xbar_demux (
		.clk                (clk_clk),                           //       clk.clk
		.reset              (rst_controller_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_src_ready),               //      sink.ready
		.sink_channel       (id_router_src_channel),             //          .channel
		.sink_data          (id_router_src_data),                //          .data
		.sink_startofpacket (id_router_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_src1_endofpacket)    //          .endofpacket
	);

	nios_system_rsp_xbar_demux_001 rsp_xbar_demux_001 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_001_src_ready),               //      sink.ready
		.sink_channel       (id_router_001_src_channel),             //          .channel
		.sink_data          (id_router_001_src_data),                //          .data
		.sink_startofpacket (id_router_001_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_001_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_001_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_001_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_001_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_001_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_001_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_001_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_001_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_001_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_001_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_001_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_001_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_001_src1_endofpacket),   //          .endofpacket
		.src2_ready         (rsp_xbar_demux_001_src2_ready),         //      src2.ready
		.src2_valid         (rsp_xbar_demux_001_src2_valid),         //          .valid
		.src2_data          (rsp_xbar_demux_001_src2_data),          //          .data
		.src2_channel       (rsp_xbar_demux_001_src2_channel),       //          .channel
		.src2_startofpacket (rsp_xbar_demux_001_src2_startofpacket), //          .startofpacket
		.src2_endofpacket   (rsp_xbar_demux_001_src2_endofpacket),   //          .endofpacket
		.src3_ready         (rsp_xbar_demux_001_src3_ready),         //      src3.ready
		.src3_valid         (rsp_xbar_demux_001_src3_valid),         //          .valid
		.src3_data          (rsp_xbar_demux_001_src3_data),          //          .data
		.src3_channel       (rsp_xbar_demux_001_src3_channel),       //          .channel
		.src3_startofpacket (rsp_xbar_demux_001_src3_startofpacket), //          .startofpacket
		.src3_endofpacket   (rsp_xbar_demux_001_src3_endofpacket)    //          .endofpacket
	);

	nios_system_cmd_xbar_demux_004 rsp_xbar_demux_002 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_002_src_ready),               //      sink.ready
		.sink_channel       (id_router_002_src_channel),             //          .channel
		.sink_data          (id_router_002_src_data),                //          .data
		.sink_startofpacket (id_router_002_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_002_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_002_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_002_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_002_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_002_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_002_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_002_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_002_src0_endofpacket)    //          .endofpacket
	);

	nios_system_rsp_xbar_demux rsp_xbar_demux_003 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_003_src_ready),               //      sink.ready
		.sink_channel       (id_router_003_src_channel),             //          .channel
		.sink_data          (id_router_003_src_data),                //          .data
		.sink_startofpacket (id_router_003_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_003_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_003_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_003_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_003_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_003_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_003_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_003_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_003_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_003_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_003_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_003_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_003_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_003_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_003_src1_endofpacket)    //          .endofpacket
	);

	nios_system_cmd_xbar_demux_004 rsp_xbar_demux_004 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_004_src_ready),               //      sink.ready
		.sink_channel       (id_router_004_src_channel),             //          .channel
		.sink_data          (id_router_004_src_data),                //          .data
		.sink_startofpacket (id_router_004_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_004_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_004_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_004_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_004_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_004_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_004_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_004_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_004_src0_endofpacket)    //          .endofpacket
	);

	nios_system_cmd_xbar_demux_004 rsp_xbar_demux_005 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_002_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_005_src_ready),               //      sink.ready
		.sink_channel       (id_router_005_src_channel),             //          .channel
		.sink_data          (id_router_005_src_data),                //          .data
		.sink_startofpacket (id_router_005_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_005_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_005_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_005_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_005_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_005_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_005_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_005_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_005_src0_endofpacket)    //          .endofpacket
	);

	nios_system_cmd_xbar_demux_004 rsp_xbar_demux_006 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_002_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_006_src_ready),               //      sink.ready
		.sink_channel       (id_router_006_src_channel),             //          .channel
		.sink_data          (id_router_006_src_data),                //          .data
		.sink_startofpacket (id_router_006_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_006_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_006_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_006_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_006_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_006_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_006_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_006_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_006_src0_endofpacket)    //          .endofpacket
	);

	nios_system_cmd_xbar_demux_004 rsp_xbar_demux_007 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_007_src_ready),               //      sink.ready
		.sink_channel       (id_router_007_src_channel),             //          .channel
		.sink_data          (id_router_007_src_data),                //          .data
		.sink_startofpacket (id_router_007_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_007_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_007_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_007_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_007_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_007_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_007_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_007_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_007_src0_endofpacket)    //          .endofpacket
	);

	nios_system_rsp_xbar_demux rsp_xbar_demux_008 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_008_src_ready),               //      sink.ready
		.sink_channel       (id_router_008_src_channel),             //          .channel
		.sink_data          (id_router_008_src_data),                //          .data
		.sink_startofpacket (id_router_008_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_008_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_008_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_008_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_008_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_008_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_008_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_008_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_008_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_008_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_008_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_008_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_008_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_008_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_008_src1_endofpacket)    //          .endofpacket
	);

	nios_system_rsp_xbar_demux rsp_xbar_demux_009 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_009_src_ready),               //      sink.ready
		.sink_channel       (id_router_009_src_channel),             //          .channel
		.sink_data          (id_router_009_src_data),                //          .data
		.sink_startofpacket (id_router_009_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_009_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_009_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_009_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_009_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_009_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_009_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_009_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_009_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_009_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_009_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_009_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_009_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_009_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_009_src1_endofpacket)    //          .endofpacket
	);

	nios_system_cmd_xbar_demux_004 rsp_xbar_demux_010 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_002_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_010_src_ready),               //      sink.ready
		.sink_channel       (id_router_010_src_channel),             //          .channel
		.sink_data          (id_router_010_src_data),                //          .data
		.sink_startofpacket (id_router_010_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_010_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_010_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_010_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_010_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_010_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_010_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_010_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_010_src0_endofpacket)    //          .endofpacket
	);

	nios_system_cmd_xbar_demux_004 rsp_xbar_demux_011 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_011_src_ready),               //      sink.ready
		.sink_channel       (id_router_011_src_channel),             //          .channel
		.sink_data          (id_router_011_src_data),                //          .data
		.sink_startofpacket (id_router_011_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_011_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_011_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_011_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_011_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_011_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_011_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_011_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_011_src0_endofpacket)    //          .endofpacket
	);

	nios_system_rsp_xbar_mux rsp_xbar_mux (
		.clk                 (clk_clk),                               //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (rsp_xbar_mux_src_ready),                //       src.ready
		.src_valid           (rsp_xbar_mux_src_valid),                //          .valid
		.src_data            (rsp_xbar_mux_src_data),                 //          .data
		.src_channel         (rsp_xbar_mux_src_channel),              //          .channel
		.src_startofpacket   (rsp_xbar_mux_src_startofpacket),        //          .startofpacket
		.src_endofpacket     (rsp_xbar_mux_src_endofpacket),          //          .endofpacket
		.sink0_ready         (rsp_xbar_demux_src0_ready),             //     sink0.ready
		.sink0_valid         (rsp_xbar_demux_src0_valid),             //          .valid
		.sink0_channel       (rsp_xbar_demux_src0_channel),           //          .channel
		.sink0_data          (rsp_xbar_demux_src0_data),              //          .data
		.sink0_startofpacket (rsp_xbar_demux_src0_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (rsp_xbar_demux_src0_endofpacket),       //          .endofpacket
		.sink1_ready         (rsp_xbar_demux_001_src0_ready),         //     sink1.ready
		.sink1_valid         (rsp_xbar_demux_001_src0_valid),         //          .valid
		.sink1_channel       (rsp_xbar_demux_001_src0_channel),       //          .channel
		.sink1_data          (rsp_xbar_demux_001_src0_data),          //          .data
		.sink1_startofpacket (rsp_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.sink1_endofpacket   (rsp_xbar_demux_001_src0_endofpacket)    //          .endofpacket
	);

	nios_system_rsp_xbar_mux_001 rsp_xbar_mux_001 (
		.clk                 (clk_clk),                               //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (rsp_xbar_mux_001_src_ready),            //       src.ready
		.src_valid           (rsp_xbar_mux_001_src_valid),            //          .valid
		.src_data            (rsp_xbar_mux_001_src_data),             //          .data
		.src_channel         (rsp_xbar_mux_001_src_channel),          //          .channel
		.src_startofpacket   (rsp_xbar_mux_001_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (rsp_xbar_mux_001_src_endofpacket),      //          .endofpacket
		.sink0_ready         (rsp_xbar_demux_src1_ready),             //     sink0.ready
		.sink0_valid         (rsp_xbar_demux_src1_valid),             //          .valid
		.sink0_channel       (rsp_xbar_demux_src1_channel),           //          .channel
		.sink0_data          (rsp_xbar_demux_src1_data),              //          .data
		.sink0_startofpacket (rsp_xbar_demux_src1_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (rsp_xbar_demux_src1_endofpacket),       //          .endofpacket
		.sink1_ready         (rsp_xbar_demux_001_src1_ready),         //     sink1.ready
		.sink1_valid         (rsp_xbar_demux_001_src1_valid),         //          .valid
		.sink1_channel       (rsp_xbar_demux_001_src1_channel),       //          .channel
		.sink1_data          (rsp_xbar_demux_001_src1_data),          //          .data
		.sink1_startofpacket (rsp_xbar_demux_001_src1_startofpacket), //          .startofpacket
		.sink1_endofpacket   (rsp_xbar_demux_001_src1_endofpacket),   //          .endofpacket
		.sink2_ready         (rsp_xbar_demux_002_src0_ready),         //     sink2.ready
		.sink2_valid         (rsp_xbar_demux_002_src0_valid),         //          .valid
		.sink2_channel       (rsp_xbar_demux_002_src0_channel),       //          .channel
		.sink2_data          (rsp_xbar_demux_002_src0_data),          //          .data
		.sink2_startofpacket (rsp_xbar_demux_002_src0_startofpacket), //          .startofpacket
		.sink2_endofpacket   (rsp_xbar_demux_002_src0_endofpacket),   //          .endofpacket
		.sink3_ready         (rsp_xbar_demux_003_src0_ready),         //     sink3.ready
		.sink3_valid         (rsp_xbar_demux_003_src0_valid),         //          .valid
		.sink3_channel       (rsp_xbar_demux_003_src0_channel),       //          .channel
		.sink3_data          (rsp_xbar_demux_003_src0_data),          //          .data
		.sink3_startofpacket (rsp_xbar_demux_003_src0_startofpacket), //          .startofpacket
		.sink3_endofpacket   (rsp_xbar_demux_003_src0_endofpacket),   //          .endofpacket
		.sink4_ready         (rsp_xbar_demux_004_src0_ready),         //     sink4.ready
		.sink4_valid         (rsp_xbar_demux_004_src0_valid),         //          .valid
		.sink4_channel       (rsp_xbar_demux_004_src0_channel),       //          .channel
		.sink4_data          (rsp_xbar_demux_004_src0_data),          //          .data
		.sink4_startofpacket (rsp_xbar_demux_004_src0_startofpacket), //          .startofpacket
		.sink4_endofpacket   (rsp_xbar_demux_004_src0_endofpacket),   //          .endofpacket
		.sink5_ready         (rsp_xbar_demux_005_src0_ready),         //     sink5.ready
		.sink5_valid         (rsp_xbar_demux_005_src0_valid),         //          .valid
		.sink5_channel       (rsp_xbar_demux_005_src0_channel),       //          .channel
		.sink5_data          (rsp_xbar_demux_005_src0_data),          //          .data
		.sink5_startofpacket (rsp_xbar_demux_005_src0_startofpacket), //          .startofpacket
		.sink5_endofpacket   (rsp_xbar_demux_005_src0_endofpacket),   //          .endofpacket
		.sink6_ready         (rsp_xbar_demux_006_src0_ready),         //     sink6.ready
		.sink6_valid         (rsp_xbar_demux_006_src0_valid),         //          .valid
		.sink6_channel       (rsp_xbar_demux_006_src0_channel),       //          .channel
		.sink6_data          (rsp_xbar_demux_006_src0_data),          //          .data
		.sink6_startofpacket (rsp_xbar_demux_006_src0_startofpacket), //          .startofpacket
		.sink6_endofpacket   (rsp_xbar_demux_006_src0_endofpacket),   //          .endofpacket
		.sink7_ready         (rsp_xbar_demux_007_src0_ready),         //     sink7.ready
		.sink7_valid         (rsp_xbar_demux_007_src0_valid),         //          .valid
		.sink7_channel       (rsp_xbar_demux_007_src0_channel),       //          .channel
		.sink7_data          (rsp_xbar_demux_007_src0_data),          //          .data
		.sink7_startofpacket (rsp_xbar_demux_007_src0_startofpacket), //          .startofpacket
		.sink7_endofpacket   (rsp_xbar_demux_007_src0_endofpacket)    //          .endofpacket
	);

	nios_system_rsp_xbar_mux_002 rsp_xbar_mux_002 (
		.clk                 (clk_clk),                               //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (rsp_xbar_mux_002_src_ready),            //       src.ready
		.src_valid           (rsp_xbar_mux_002_src_valid),            //          .valid
		.src_data            (rsp_xbar_mux_002_src_data),             //          .data
		.src_channel         (rsp_xbar_mux_002_src_channel),          //          .channel
		.src_startofpacket   (rsp_xbar_mux_002_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (rsp_xbar_mux_002_src_endofpacket),      //          .endofpacket
		.sink0_ready         (rsp_xbar_demux_003_src1_ready),         //     sink0.ready
		.sink0_valid         (rsp_xbar_demux_003_src1_valid),         //          .valid
		.sink0_channel       (rsp_xbar_demux_003_src1_channel),       //          .channel
		.sink0_data          (rsp_xbar_demux_003_src1_data),          //          .data
		.sink0_startofpacket (rsp_xbar_demux_003_src1_startofpacket), //          .startofpacket
		.sink0_endofpacket   (rsp_xbar_demux_003_src1_endofpacket),   //          .endofpacket
		.sink1_ready         (rsp_xbar_demux_008_src0_ready),         //     sink1.ready
		.sink1_valid         (rsp_xbar_demux_008_src0_valid),         //          .valid
		.sink1_channel       (rsp_xbar_demux_008_src0_channel),       //          .channel
		.sink1_data          (rsp_xbar_demux_008_src0_data),          //          .data
		.sink1_startofpacket (rsp_xbar_demux_008_src0_startofpacket), //          .startofpacket
		.sink1_endofpacket   (rsp_xbar_demux_008_src0_endofpacket),   //          .endofpacket
		.sink2_ready         (rsp_xbar_demux_009_src0_ready),         //     sink2.ready
		.sink2_valid         (rsp_xbar_demux_009_src0_valid),         //          .valid
		.sink2_channel       (rsp_xbar_demux_009_src0_channel),       //          .channel
		.sink2_data          (rsp_xbar_demux_009_src0_data),          //          .data
		.sink2_startofpacket (rsp_xbar_demux_009_src0_startofpacket), //          .startofpacket
		.sink2_endofpacket   (rsp_xbar_demux_009_src0_endofpacket),   //          .endofpacket
		.sink3_ready         (rsp_xbar_demux_010_src0_ready),         //     sink3.ready
		.sink3_valid         (rsp_xbar_demux_010_src0_valid),         //          .valid
		.sink3_channel       (rsp_xbar_demux_010_src0_channel),       //          .channel
		.sink3_data          (rsp_xbar_demux_010_src0_data),          //          .data
		.sink3_startofpacket (rsp_xbar_demux_010_src0_startofpacket), //          .startofpacket
		.sink3_endofpacket   (rsp_xbar_demux_010_src0_endofpacket),   //          .endofpacket
		.sink4_ready         (rsp_xbar_demux_011_src0_ready),         //     sink4.ready
		.sink4_valid         (rsp_xbar_demux_011_src0_valid),         //          .valid
		.sink4_channel       (rsp_xbar_demux_011_src0_channel),       //          .channel
		.sink4_data          (rsp_xbar_demux_011_src0_data),          //          .data
		.sink4_startofpacket (rsp_xbar_demux_011_src0_startofpacket), //          .startofpacket
		.sink4_endofpacket   (rsp_xbar_demux_011_src0_endofpacket)    //          .endofpacket
	);

	nios_system_rsp_xbar_mux rsp_xbar_mux_003 (
		.clk                 (clk_clk),                               //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (rsp_xbar_mux_003_src_ready),            //       src.ready
		.src_valid           (rsp_xbar_mux_003_src_valid),            //          .valid
		.src_data            (rsp_xbar_mux_003_src_data),             //          .data
		.src_channel         (rsp_xbar_mux_003_src_channel),          //          .channel
		.src_startofpacket   (rsp_xbar_mux_003_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (rsp_xbar_mux_003_src_endofpacket),      //          .endofpacket
		.sink0_ready         (rsp_xbar_demux_008_src1_ready),         //     sink0.ready
		.sink0_valid         (rsp_xbar_demux_008_src1_valid),         //          .valid
		.sink0_channel       (rsp_xbar_demux_008_src1_channel),       //          .channel
		.sink0_data          (rsp_xbar_demux_008_src1_data),          //          .data
		.sink0_startofpacket (rsp_xbar_demux_008_src1_startofpacket), //          .startofpacket
		.sink0_endofpacket   (rsp_xbar_demux_008_src1_endofpacket),   //          .endofpacket
		.sink1_ready         (rsp_xbar_demux_009_src1_ready),         //     sink1.ready
		.sink1_valid         (rsp_xbar_demux_009_src1_valid),         //          .valid
		.sink1_channel       (rsp_xbar_demux_009_src1_channel),       //          .channel
		.sink1_data          (rsp_xbar_demux_009_src1_data),          //          .data
		.sink1_startofpacket (rsp_xbar_demux_009_src1_startofpacket), //          .startofpacket
		.sink1_endofpacket   (rsp_xbar_demux_009_src1_endofpacket)    //          .endofpacket
	);

	nios_system_cmd_xbar_demux_006 cmd_xbar_demux_006 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (addr_router_006_src_ready),             //      sink.ready
		.sink_channel       (addr_router_006_src_channel),           //          .channel
		.sink_data          (addr_router_006_src_data),              //          .data
		.sink_startofpacket (addr_router_006_src_startofpacket),     //          .startofpacket
		.sink_endofpacket   (addr_router_006_src_endofpacket),       //          .endofpacket
		.sink_valid         (addr_router_006_src_valid),             //          .valid
		.src0_ready         (cmd_xbar_demux_006_src0_ready),         //      src0.ready
		.src0_valid         (cmd_xbar_demux_006_src0_valid),         //          .valid
		.src0_data          (cmd_xbar_demux_006_src0_data),          //          .data
		.src0_channel       (cmd_xbar_demux_006_src0_channel),       //          .channel
		.src0_startofpacket (cmd_xbar_demux_006_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_006_src0_endofpacket)    //          .endofpacket
	);

	nios_system_cmd_xbar_demux_006 rsp_xbar_demux_012 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_012_src_ready),               //      sink.ready
		.sink_channel       (id_router_012_src_channel),             //          .channel
		.sink_data          (id_router_012_src_data),                //          .data
		.sink_startofpacket (id_router_012_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_012_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_012_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_012_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_012_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_012_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_012_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_012_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_012_src0_endofpacket)    //          .endofpacket
	);

	nios_system_cmd_xbar_demux_006 cmd_xbar_demux_007 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (addr_router_007_src_ready),             //      sink.ready
		.sink_channel       (addr_router_007_src_channel),           //          .channel
		.sink_data          (addr_router_007_src_data),              //          .data
		.sink_startofpacket (addr_router_007_src_startofpacket),     //          .startofpacket
		.sink_endofpacket   (addr_router_007_src_endofpacket),       //          .endofpacket
		.sink_valid         (addr_router_007_src_valid),             //          .valid
		.src0_ready         (cmd_xbar_demux_007_src0_ready),         //      src0.ready
		.src0_valid         (cmd_xbar_demux_007_src0_valid),         //          .valid
		.src0_data          (cmd_xbar_demux_007_src0_data),          //          .data
		.src0_channel       (cmd_xbar_demux_007_src0_channel),       //          .channel
		.src0_startofpacket (cmd_xbar_demux_007_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_007_src0_endofpacket)    //          .endofpacket
	);

	nios_system_cmd_xbar_demux_006 rsp_xbar_demux_013 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_013_src_ready),               //      sink.ready
		.sink_channel       (id_router_013_src_channel),             //          .channel
		.sink_data          (id_router_013_src_data),                //          .data
		.sink_startofpacket (id_router_013_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_013_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_013_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_013_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_013_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_013_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_013_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_013_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_013_src0_endofpacket)    //          .endofpacket
	);

	nios_system_irq_mapper irq_mapper (
		.clk           (clk_clk),                        //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),       // receiver2.irq
		.receiver3_irq (irq_mapper_receiver3_irq),       // receiver3.irq
		.sender_irq    (com_nios_d_irq_irq)              //    sender.irq
	);

	nios_system_irq_mapper_001 irq_mapper_001 (
		.clk           (clk_clk),                        //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_001_receiver0_irq),   // receiver0.irq
		.sender_irq    (carcontrol_nios_d_irq_irq)       //    sender.irq
	);

endmodule
